module MemInst(
    input [31:0] pc,          // endereço de instrução (program counter)
    output reg [31:0] out_inst,   // saída de instrução (16 bits)
    input clock,
    input stall
);


    // Memória de instruções (256 posições, 8 bits cada)
    reg [7:0] inst [0:255];

    // Inicialização das memórias

    initial begin //addi,add,sub,jalr e jal(nsalva pc atual, não anterior), sll, or, sra, srl, blt, auipc, lui, lw, sw
    //inst[0] = 32'b00000000-0001_0000-0_000_0001-0_0010011; //addi 2 0 1
    //inst[1] = 32'b0000000_00010_00010_000_00001_0110011; //add 1 0 2
    //inst[2] = 32'b0000000_00001_00000_010_00100_0100011; //sw valor 1 --> 4
    //inst[3] = 32'b000000000100_00000_010_00100_0000011; //lw valor 4 --> 4
    //inst[2] = 32'b00000000000000000010_11111_0010111; //auipc pc + 2
    //inst[2] = 32'b10000000000000000000_11111_0110111; //lui 1 no mais significativo
    //inst[2] = 32'b0000000_00001_00010_100_10100_1100011; //blt pc+10 1 2
    //inst[3] = 32'b0000000_00010_00010_100_10100_1100011; //blt pc+10 1 1
    //inst[2] = 32'b0100000_00010_00001_100_00011_0110011; //sra 3 2 1
    //inst[3] = 32'b0100000_00010_00001_110_00011_0110011; // or 3 2 1
    //inst[4] = 32'b0100000_00010_00001_001_00011_0110011; // sll 3 2 1
    //inst[3] = 32'b0100000_00010_00001_101_00011_0110011; // srl 3 2 1
    //inst[7] = 32'b0100000_00010_00001_011_00011_0110011; //sub 3 2 1
    //inst[3] = 32'b000000001010_00001_000_11111_1100111; //jalr 2 + 10
    //inst[4] = 32'b00000000000000000001_11111_1101111; //jal 1 11111
    //inst[4] = 32'b00000000000000000001_00111_0010111; //aui pc +1, 7
    //inst[5] = 32'b11000000000000000001_11111_0110111; //lui 11...00001 11


    //addi 2 0 4
    /*
    inst[0] = 8'b00000000;
    inst[1] = 8'b01000000;
    inst[2] = 8'b00000001;
    inst[3] = 8'b00010011;

    inst[4] = 8'b00000000;
    inst[5] = 8'b00000000;
    inst[6] = 8'b00000000;
    inst[7] = 8'b00000000;

    inst[8] = 8'b00000000;
    inst[9] = 8'b00000000;
    inst[10] = 8'b00000000;
    inst[11] = 8'b00000000;

    inst[12] = 8'b00000000;
    inst[13] = 8'b00000000;
    inst[14] = 8'b00000000;
    inst[15] = 8'b00000000;


    //jalr 2 + 12
    inst[16] = 8'b00000000;
    inst[17] = 8'b1100_0001;
    inst[18] = 8'b0_000_1111;
    inst[19] = 8'b1_1100111;

    inst[20] = 8'b00000000;
    inst[21] = 8'b00000000;
    inst[22] = 8'b00000000;
    inst[23] = 8'b00000000;

    inst[24] = 8'b00000000;
    inst[25] = 8'b00000000;
    inst[26] = 8'b00000000;
    inst[27] = 8'b00000000;

    inst[28] = 8'b00000000;
    inst[29] = 8'b00000000;
    inst[30] = 8'b00000000;
    inst[31] = 8'b00000000;
    */

    // jal test
inst[0] = 8'b11111000;
inst[1] = 8'b00000000;
inst[2] = 8'b00011111;
inst[3] = 8'b11101111;
// addi 2 0 1
inst[4] = 8'b00000000;
inst[5] = 8'b00010000;
inst[6] = 8'b00000001;
inst[7] = 8'b00010011;
// addi 3 0 2
inst[8] = 8'b00000000;
inst[9] = 8'b00100000;
inst[10] = 8'b00000001;
inst[11] = 8'b10010011;
// add 1 3 2
inst[12] = 8'b00000000;
inst[13] = 8'b00110001;
inst[14] = 8'b00000000;
inst[15] = 8'b10110011;
// add 4 3 2
inst[16] = 8'b00000000;
inst[17] = 8'b00110001;
inst[18] = 8'b00000010;
inst[19] = 8'b00110011;
// add 5 3 2
inst[20] = 8'b00000000;
inst[21] = 8'b00110001;
inst[22] = 8'b00000010;
inst[23] = 8'b10110011;
    /*
    //jal 32 11111
    inst[16] = 8'b00000000;
    inst[17] = 8'b00000010;
    inst[18] = 8'b0000_1111;
    inst[19] = 8'b1_1101111;

    inst[20] = 8'b00000000;
    inst[21] = 8'b00000000;
    inst[22] = 8'b00000000;
    inst[23] = 8'b00000000;

    inst[24] = 8'b00000000;
    inst[25] = 8'b00000000;
    inst[26] = 8'b00000000;
    inst[27] = 8'b00000000;

    inst[28] = 8'b00000000;
    inst[29] = 8'b00000000;
    inst[30] = 8'b00000000;
    inst[31] = 8'b00000000;
    */


    /*
    //addi 2 0 1
    inst[0] = 8'b00000000;
    inst[1] = 8'b00010000;
    inst[2] = 8'b00000001;
    inst[3] = 8'b00010011;

    inst[4] = 8'b00000000;
    inst[5] = 8'b00000000;
    inst[6] = 8'b00000000;
    inst[7] = 8'b00000000;

    inst[8] = 8'b00000000;
    inst[9] = 8'b00000000;
    inst[10] = 8'b00000000;
    inst[11] = 8'b00000000;

    inst[12] = 8'b00000000;
    inst[13] = 8'b00000000;
    inst[14] = 8'b00000000;
    inst[15] = 8'b00000000;

    //add 6 2 1
    inst[16] = 8'b00000000;
    inst[17] = 8'b00010001;
    inst[18] = 8'b00000011;
    inst[19] = 8'b00010011;

    inst[20] = 8'b00000000;
    inst[21] = 8'b00000000;
    inst[22] = 8'b00000000;
    inst[23] = 8'b00000000;

    inst[24] = 8'b00000000;
    inst[25] = 8'b00000000;
    inst[26] = 8'b00000000;
    inst[27] = 8'b00000000;

    inst[28] = 8'b00000000;
    inst[29] = 8'b00000000;
    inst[30] = 8'b00000000;
    inst[31] = 8'b00000000;

    //sub 3 2 1
    inst[32] = 8'b0100000_0;
    inst[33] = 8'b0010_0000;
    inst[34] = 8'b1_011_0001;
    inst[35] = 8'b1_0110011;

    inst[36] = 8'b00000000;
    inst[37] = 8'b00000000;
    inst[38] = 8'b00000000;
    inst[39] = 8'b00000000;

    inst[40] = 8'b00000000;
    inst[41] = 8'b00000000;
    inst[42] = 8'b00000000;
    inst[43] = 8'b00000000;

    inst[44] = 8'b00000000;
    inst[45] = 8'b00000000;
    inst[46] = 8'b00000000;
    inst[47] = 8'b00000000;

    //sw valor 3 --> 4
    inst[48] = 8'b0000000_0;
    inst[49] = 8'b0011_0000;
    inst[50] = 8'b0_010_0010;
    inst[51] = 8'b0_0100011;

    inst[52] = 8'b00000000;
    inst[53] = 8'b00000000;
    inst[54] = 8'b00000000;
    inst[55] = 8'b00000000;

    inst[56] = 8'b00000000;
    inst[57] = 8'b00000000;
    inst[58] = 8'b00000000;
    inst[59] = 8'b00000000;

    inst[60] = 8'b00000000;
    inst[61] = 8'b00000000;
    inst[62] = 8'b00000000;
    inst[63] = 8'b00000000;

    //lw valor 4 --> 4
    inst[64] = 8'b00000000;
    inst[65] = 8'b0100_0000;
    inst[66] = 8'b0_010_0010;
    inst[67] = 8'b0_0000011;

    inst[68] = 8'b00000000;
    inst[69] = 8'b00000000;
    inst[70] = 8'b00000000;
    inst[71] = 8'b00000000;

    inst[72] = 8'b00000000;
    inst[73] = 8'b00000000;
    inst[74] = 8'b00000000;
    inst[75] = 8'b00000000;

    inst[76] = 8'b00000000;
    inst[77] = 8'b00000000;
    inst[78] = 8'b00000000;
    inst[79] = 8'b00000000;

    //auipc pc + 2 --> 31
    inst[80] = 8'b00000000;
    inst[81] = 8'b00000000;
    inst[82] = 8'b0010_1111;
    inst[83] = 8'b1_0010111;

    inst[84] = 8'b00000000;
    inst[85] = 8'b00000000;
    inst[86] = 8'b00000000;
    inst[87] = 8'b00000000;

    inst[88] = 8'b00000000;
    inst[89] = 8'b00000000;
    inst[90] = 8'b00000000;
    inst[91] = 8'b00000000;

    inst[92] = 8'b00000000;
    inst[93] = 8'b00000000;
    inst[94] = 8'b00000000;
    inst[95] = 8'b00000000;

    //lui 1 no mais significativo
    inst[96] = 8'b10000000;
    inst[97] = 8'b00000000;
    inst[98] = 8'b0000_1111;
    inst[99] = 8'b1_0110111;

    inst[100] = 8'b00000000;
    inst[101] = 8'b00000000;
    inst[102] = 8'b00000000;
    inst[103] = 8'b00000000;

    inst[104] = 8'b00000000;
    inst[105] = 8'b00000000;
    inst[106] = 8'b00000000;
    inst[107] = 8'b00000000;

    inst[108] = 8'b00000000;
    inst[109] = 8'b00000000;
    inst[110] = 8'b00000000;
    inst[111] = 8'b00000000;

    //blt pc+10 1 2
    inst[112] = 8'b0000000_0;
    inst[113] = 8'b0001_0001;
    inst[114] = 8'b0_100_1000;
    inst[115] = 8'b0_1100011;

    inst[116] = 8'b00000000;
    inst[117] = 8'b00000000;
    inst[118] = 8'b00000000;
    inst[119] = 8'b00000000;

    inst[120] = 8'b00000000;
    inst[121] = 8'b00000000;
    inst[122] = 8'b00000000;
    inst[123] = 8'b00000000;

    inst[124] = 8'b00000000;
    inst[125] = 8'b00000000;
    inst[126] = 8'b00000000;
    inst[127] = 8'b00000000;

    //blt pc+10 1 1
    inst[128] = 8'b0000000_0;
    inst[129] = 8'b001_00000_;
    inst[130] = 8'b010_01000;
    inst[131] = 8'b0_1100011;

    inst[132] = 8'b00000000;
    inst[133] = 8'b00000000;
    inst[134] = 8'b00000000;
    inst[135]= 8'b00000000;

    inst[136] = 8'b00000000;
    inst[137] = 8'b00000000;
    inst[138] = 8'b00000000;
    inst[139] = 8'b00000000;

    inst[140] = 8'b00000000;
    inst[141] = 8'b00000000;
    inst[142] = 8'b00000000;
    inst[143] = 8'b00000000;
    */
        // ... (inicialize o restante das posições com 0)

        // Instruções já fornecidas

        // ... (inicialize o restante das instruções com 0)
    end

    always @(posedge clock, posedge stall)

    begin
    if (stall)
        begin
        out_inst <= 32'b0;
        end
    else
        out_inst <= {inst[pc], inst[pc+1], inst[pc+2], inst[pc+3]};     // Saída de instrução
    end

endmodule
