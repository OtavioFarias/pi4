module MemDat(
    input [31:0] value,       // valor de entrada (8 bits)
    input esc_mem,           // sinal de controle para escrita em memória
    input read_mem,
    input [31:0] dst_mem,     // endereço de destino para escrita
    output [31:0] out_dat,  // saída de dados (8 bits)
    input clock
);
//colocar readMem
    // Memória de dados (256 posições, 8 bits cada)
    reg [7:0] dat [0:4095];

    // Inicialização das memórias
    initial begin

dat[0] = 8'b00000000;
dat[1] = 8'b00000000;
dat[2] = 8'b00000000;
dat[3] = 8'b00000001;

dat[4] = 8'b00000000;
dat[5] = 8'b00000000;
dat[6] = 8'b00000000;
dat[7] = 8'b00000010;

dat[8] = 8'b00000000;
dat[9] = 8'b00000000;
dat[10] = 8'b00000000;
dat[11] = 8'b00000101;

dat[12] = 8'b00000000;
dat[13] = 8'b00000000;
dat[14] = 8'b00000000;
dat[15] = 8'b00000100;

dat[16] = 8'b00000000;
dat[17] = 8'b00000000;
dat[18] = 8'b00000000;
dat[19] = 8'b00000000;
dat[20] = 8'b00000000;
dat[21] = 8'b00000000;
dat[22] = 8'b00000000;
dat[23] = 8'b00000000;
dat[24] = 8'b00000000;
dat[25] = 8'b00000000;
dat[26] = 8'b00000000;
dat[27] = 8'b00000000;
dat[28] = 8'b00000000;
dat[29] = 8'b00000000;
dat[30] = 8'b00000000;
dat[31] = 8'b00000000;
dat[32] = 8'b00000000;
dat[33] = 8'b00000000;
dat[34] = 8'b00000000;
dat[35] = 8'b00000000;
dat[36] = 8'b00000000;
dat[37] = 8'b00000000;
dat[38] = 8'b00000000;
dat[39] = 8'b00000000;
dat[40] = 8'b00000000;
dat[41] = 8'b00000000;
dat[42] = 8'b00000000;
dat[43] = 8'b00000000;
dat[44] = 8'b00000000;
dat[45] = 8'b00000000;
dat[46] = 8'b00000000;
dat[47] = 8'b00000000;
dat[48] = 8'b00000000;
dat[49] = 8'b00000000;
dat[50] = 8'b00000000;
dat[51] = 8'b00000000;
dat[52] = 8'b00000000;
dat[53] = 8'b00000000;
dat[54] = 8'b00000000;
dat[55] = 8'b00000000;
dat[56] = 8'b00000000;
dat[57] = 8'b00000000;
dat[58] = 8'b00000000;
dat[59] = 8'b00000000;
dat[60] = 8'b00000000;
dat[61] = 8'b00000000;
dat[62] = 8'b00000000;
dat[63] = 8'b00000000;
dat[64] = 8'b00000000;
dat[65] = 8'b00000000;
dat[66] = 8'b00000000;
dat[67] = 8'b00000000;
dat[68] = 8'b00000000;
dat[69] = 8'b00000000;
dat[70] = 8'b00000000;
dat[71] = 8'b00000000;
dat[72] = 8'b00000000;
dat[73] = 8'b00000000;
dat[74] = 8'b00000000;
dat[75] = 8'b00000000;
dat[76] = 8'b00000000;
dat[77] = 8'b00000000;
dat[78] = 8'b00000000;
dat[79] = 8'b00000000;
dat[80] = 8'b00000000;
dat[81] = 8'b00000000;
dat[82] = 8'b00000000;
dat[83] = 8'b00000000;
dat[84] = 8'b00000000;
dat[85] = 8'b00000000;
dat[86] = 8'b00000000;
dat[87] = 8'b00000000;
dat[88] = 8'b00000000;
dat[89] = 8'b00000000;
dat[90] = 8'b00000000;
dat[91] = 8'b00000000;
dat[92] = 8'b00000000;
dat[93] = 8'b00000000;
dat[94] = 8'b00000000;
dat[95] = 8'b00000000;
dat[96] = 8'b00000000;
dat[97] = 8'b00000000;
dat[98] = 8'b00000000;
dat[99] = 8'b00000000;
dat[100] = 8'b00000000;
dat[101] = 8'b00000000;
dat[102] = 8'b00000000;
dat[103] = 8'b00000000;
dat[104] = 8'b00000000;
dat[105] = 8'b00000000;
dat[106] = 8'b00000000;
dat[107] = 8'b00000000;
dat[108] = 8'b00000000;
dat[109] = 8'b00000000;
dat[110] = 8'b00000000;
dat[111] = 8'b00000000;
dat[112] = 8'b00000000;
dat[113] = 8'b00000000;
dat[114] = 8'b00000000;
dat[115] = 8'b00000000;
dat[116] = 8'b00000000;
dat[117] = 8'b00000000;
dat[118] = 8'b00000000;
dat[119] = 8'b00000000;
dat[120] = 8'b00000000;
dat[121] = 8'b00000000;
dat[122] = 8'b00000000;
dat[123] = 8'b00000000;
dat[124] = 8'b00000000;
dat[125] = 8'b00000000;
dat[126] = 8'b00000000;
dat[127] = 8'b00000000;
dat[128] = 8'b00000000;
dat[129] = 8'b00000000;
dat[130] = 8'b00000000;
dat[131] = 8'b00000000;
dat[132] = 8'b00000000;
dat[133] = 8'b00000000;
dat[134] = 8'b00000000;
dat[135] = 8'b00000000;
dat[136] = 8'b00000000;
dat[137] = 8'b00000000;
dat[138] = 8'b00000000;
dat[139] = 8'b00000000;
dat[140] = 8'b00000000;
dat[141] = 8'b00000000;
dat[142] = 8'b00000000;
dat[143] = 8'b00000000;
dat[144] = 8'b00000000;
dat[145] = 8'b00000000;
dat[146] = 8'b00000000;
dat[147] = 8'b00000000;
dat[148] = 8'b00000000;
dat[149] = 8'b00000000;
dat[150] = 8'b00000000;
dat[151] = 8'b00000000;
dat[152] = 8'b00000000;
dat[153] = 8'b00000000;
dat[154] = 8'b00000000;
dat[155] = 8'b00000000;
dat[156] = 8'b00000000;
dat[157] = 8'b00000000;
dat[158] = 8'b00000000;
dat[159] = 8'b00000000;
dat[160] = 8'b00000000;
dat[161] = 8'b00000000;
dat[162] = 8'b00000000;
dat[163] = 8'b00000000;
dat[164] = 8'b00000000;
dat[165] = 8'b00000000;
dat[166] = 8'b00000000;
dat[167] = 8'b00000000;
dat[168] = 8'b00000000;
dat[169] = 8'b00000000;
dat[170] = 8'b00000000;
dat[171] = 8'b00000000;
dat[172] = 8'b00000000;
dat[173] = 8'b00000000;
dat[174] = 8'b00000000;
dat[175] = 8'b00000000;
dat[176] = 8'b00000000;
dat[177] = 8'b00000000;
dat[178] = 8'b00000000;
dat[179] = 8'b00000000;
dat[180] = 8'b00000000;
dat[181] = 8'b00000000;
dat[182] = 8'b00000000;
dat[183] = 8'b00000000;
dat[184] = 8'b00000000;
dat[185] = 8'b00000000;
dat[186] = 8'b00000000;
dat[187] = 8'b00000000;
dat[188] = 8'b00000000;
dat[189] = 8'b00000000;
dat[190] = 8'b00000000;
dat[191] = 8'b00000000;
dat[192] = 8'b00000000;
dat[193] = 8'b00000000;
dat[194] = 8'b00000000;
dat[195] = 8'b00000000;
dat[196] = 8'b00000000;
dat[197] = 8'b00000000;
dat[198] = 8'b00000000;
dat[199] = 8'b00000000;
dat[200] = 8'b00000000;
dat[201] = 8'b00000000;
dat[202] = 8'b00000000;
dat[203] = 8'b00000000;
dat[204] = 8'b00000000;
dat[205] = 8'b00000000;
dat[206] = 8'b00000000;
dat[207] = 8'b00000000;
dat[208] = 8'b00000000;
dat[209] = 8'b00000000;
dat[210] = 8'b00000000;
dat[211] = 8'b00000000;
dat[212] = 8'b00000000;
dat[213] = 8'b00000000;
dat[214] = 8'b00000000;
dat[215] = 8'b00000000;
dat[216] = 8'b00000000;
dat[217] = 8'b00000000;
dat[218] = 8'b00000000;
dat[219] = 8'b00000000;
dat[220] = 8'b00000000;
dat[221] = 8'b00000000;
dat[222] = 8'b00000000;
dat[223] = 8'b00000000;
dat[224] = 8'b00000000;
dat[225] = 8'b00000000;
dat[226] = 8'b00000000;
dat[227] = 8'b00000000;
dat[228] = 8'b00000000;
dat[229] = 8'b00000000;
dat[230] = 8'b00000000;
dat[231] = 8'b00000000;
dat[232] = 8'b00000000;
dat[233] = 8'b00000000;
dat[234] = 8'b00000000;
dat[235] = 8'b00000000;
dat[236] = 8'b00000000;
dat[237] = 8'b00000000;
dat[238] = 8'b00000000;
dat[239] = 8'b00000000;
dat[240] = 8'b00000000;
dat[241] = 8'b00000000;
dat[242] = 8'b00000000;
dat[243] = 8'b00000000;
dat[244] = 8'b00000000;
dat[245] = 8'b00000000;
dat[246] = 8'b00000000;
dat[247] = 8'b00000000;
dat[248] = 8'b00000000;
dat[249] = 8'b00000000;
dat[250] = 8'b00000000;
dat[251] = 8'b00000000;
dat[252] = 8'b00000000;
dat[253] = 8'b00000000;
dat[254] = 8'b00000000;
dat[255] = 8'b00000000;
dat[256] = 8'b00000000;
dat[257] = 8'b00000000;
dat[258] = 8'b00000000;
dat[259] = 8'b00000000;
dat[260] = 8'b00000000;
dat[261] = 8'b00000000;
dat[262] = 8'b00000000;
dat[263] = 8'b00000000;
dat[264] = 8'b00000000;
dat[265] = 8'b00000000;
dat[266] = 8'b00000000;
dat[267] = 8'b00000000;
dat[268] = 8'b00000000;
dat[269] = 8'b00000000;
dat[270] = 8'b00000000;
dat[271] = 8'b00000000;
dat[272] = 8'b00000000;
dat[273] = 8'b00000000;
dat[274] = 8'b00000000;
dat[275] = 8'b00000000;
dat[276] = 8'b00000000;
dat[277] = 8'b00000000;
dat[278] = 8'b00000000;
dat[279] = 8'b00000000;
dat[280] = 8'b00000000;
dat[281] = 8'b00000000;
dat[282] = 8'b00000000;
dat[283] = 8'b00000000;
dat[284] = 8'b00000000;
dat[285] = 8'b00000000;
dat[286] = 8'b00000000;
dat[287] = 8'b00000000;
dat[288] = 8'b00000000;
dat[289] = 8'b00000000;
dat[290] = 8'b00000000;
dat[291] = 8'b00000000;
dat[292] = 8'b00000000;
dat[293] = 8'b00000000;
dat[294] = 8'b00000000;
dat[295] = 8'b00000000;
dat[296] = 8'b00000000;
dat[297] = 8'b00000000;
dat[298] = 8'b00000000;
dat[299] = 8'b00000000;
dat[300] = 8'b00000000;
dat[301] = 8'b00000000;
dat[302] = 8'b00000000;
dat[303] = 8'b00000000;
dat[304] = 8'b00000000;
dat[305] = 8'b00000000;
dat[306] = 8'b00000000;
dat[307] = 8'b00000000;
dat[308] = 8'b00000000;
dat[309] = 8'b00000000;
dat[310] = 8'b00000000;
dat[311] = 8'b00000000;
dat[312] = 8'b00000000;
dat[313] = 8'b00000000;
dat[314] = 8'b00000000;
dat[315] = 8'b00000000;
dat[316] = 8'b00000000;
dat[317] = 8'b00000000;
dat[318] = 8'b00000000;
dat[319] = 8'b00000000;
dat[320] = 8'b00000000;
dat[321] = 8'b00000000;
dat[322] = 8'b00000000;
dat[323] = 8'b00000000;
dat[324] = 8'b00000000;
dat[325] = 8'b00000000;
dat[326] = 8'b00000000;
dat[327] = 8'b00000000;
dat[328] = 8'b00000000;
dat[329] = 8'b00000000;
dat[330] = 8'b00000000;
dat[331] = 8'b00000000;
dat[332] = 8'b00000000;
dat[333] = 8'b00000000;
dat[334] = 8'b00000000;
dat[335] = 8'b00000000;
dat[336] = 8'b00000000;
dat[337] = 8'b00000000;
dat[338] = 8'b00000000;
dat[339] = 8'b00000000;
dat[340] = 8'b00000000;
dat[341] = 8'b00000000;
dat[342] = 8'b00000000;
dat[343] = 8'b00000000;
dat[344] = 8'b00000000;
dat[345] = 8'b00000000;
dat[346] = 8'b00000000;
dat[347] = 8'b00000000;
dat[348] = 8'b00000000;
dat[349] = 8'b00000000;
dat[350] = 8'b00000000;
dat[351] = 8'b00000000;
dat[352] = 8'b00000000;
dat[353] = 8'b00000000;
dat[354] = 8'b00000000;
dat[355] = 8'b00000000;
dat[356] = 8'b00000000;
dat[357] = 8'b00000000;
dat[358] = 8'b00000000;
dat[359] = 8'b00000000;
dat[360] = 8'b00000000;
dat[361] = 8'b00000000;
dat[362] = 8'b00000000;
dat[363] = 8'b00000000;
dat[364] = 8'b00000000;
dat[365] = 8'b00000000;
dat[366] = 8'b00000000;
dat[367] = 8'b00000000;
dat[368] = 8'b00000000;
dat[369] = 8'b00000000;
dat[370] = 8'b00000000;
dat[371] = 8'b00000000;
dat[372] = 8'b00000000;
dat[373] = 8'b00000000;
dat[374] = 8'b00000000;
dat[375] = 8'b00000000;
dat[376] = 8'b00000000;
dat[377] = 8'b00000000;
dat[378] = 8'b00000000;
dat[379] = 8'b00000000;
dat[380] = 8'b00000000;
dat[381] = 8'b00000000;
dat[382] = 8'b00000000;
dat[383] = 8'b00000000;
dat[384] = 8'b00000000;
dat[385] = 8'b00000000;
dat[386] = 8'b00000000;
dat[387] = 8'b00000000;
dat[388] = 8'b00000000;
dat[389] = 8'b00000000;
dat[390] = 8'b00000000;
dat[391] = 8'b00000000;
dat[392] = 8'b00000000;
dat[393] = 8'b00000000;
dat[394] = 8'b00000000;
dat[395] = 8'b00000000;
dat[396] = 8'b00000000;
dat[397] = 8'b00000000;
dat[398] = 8'b00000000;
dat[399] = 8'b00000000;
dat[400] = 8'b00000000;
dat[401] = 8'b00000000;
dat[402] = 8'b00000000;
dat[403] = 8'b00000000;
dat[404] = 8'b00000000;
dat[405] = 8'b00000000;
dat[406] = 8'b00000000;
dat[407] = 8'b00000000;
dat[408] = 8'b00000000;
dat[409] = 8'b00000000;
dat[410] = 8'b00000000;
dat[411] = 8'b00000000;
dat[412] = 8'b00000000;
dat[413] = 8'b00000000;
dat[414] = 8'b00000000;
dat[415] = 8'b00000000;
dat[416] = 8'b00000000;
dat[417] = 8'b00000000;
dat[418] = 8'b00000000;
dat[419] = 8'b00000000;
dat[420] = 8'b00000000;
dat[421] = 8'b00000000;
dat[422] = 8'b00000000;
dat[423] = 8'b00000000;
dat[424] = 8'b00000000;
dat[425] = 8'b00000000;
dat[426] = 8'b00000000;
dat[427] = 8'b00000000;
dat[428] = 8'b00000000;
dat[429] = 8'b00000000;
dat[430] = 8'b00000000;
dat[431] = 8'b00000000;
dat[432] = 8'b00000000;
dat[433] = 8'b00000000;
dat[434] = 8'b00000000;
dat[435] = 8'b00000000;
dat[436] = 8'b00000000;
dat[437] = 8'b00000000;
dat[438] = 8'b00000000;
dat[439] = 8'b00000000;
dat[440] = 8'b00000000;
dat[441] = 8'b00000000;
dat[442] = 8'b00000000;
dat[443] = 8'b00000000;
dat[444] = 8'b00000000;
dat[445] = 8'b00000000;
dat[446] = 8'b00000000;
dat[447] = 8'b00000000;
dat[448] = 8'b00000000;
dat[449] = 8'b00000000;
dat[450] = 8'b00000000;
dat[451] = 8'b00000000;
dat[452] = 8'b00000000;
dat[453] = 8'b00000000;
dat[454] = 8'b00000000;
dat[455] = 8'b00000000;
dat[456] = 8'b00000000;
dat[457] = 8'b00000000;
dat[458] = 8'b00000000;
dat[459] = 8'b00000000;
dat[460] = 8'b00000000;
dat[461] = 8'b00000000;
dat[462] = 8'b00000000;
dat[463] = 8'b00000000;
dat[464] = 8'b00000000;
dat[465] = 8'b00000000;
dat[466] = 8'b00000000;
dat[467] = 8'b00000000;
dat[468] = 8'b00000000;
dat[469] = 8'b00000000;
dat[470] = 8'b00000000;
dat[471] = 8'b00000000;
dat[472] = 8'b00000000;
dat[473] = 8'b00000000;
dat[474] = 8'b00000000;
dat[475] = 8'b00000000;
dat[476] = 8'b00000000;
dat[477] = 8'b00000000;
dat[478] = 8'b00000000;
dat[479] = 8'b00000000;
dat[480] = 8'b00000000;
dat[481] = 8'b00000000;
dat[482] = 8'b00000000;
dat[483] = 8'b00000000;
dat[484] = 8'b00000000;
dat[485] = 8'b00000000;
dat[486] = 8'b00000000;
dat[487] = 8'b00000000;
dat[488] = 8'b00000000;
dat[489] = 8'b00000000;
dat[490] = 8'b00000000;
dat[491] = 8'b00000000;
dat[492] = 8'b00000000;
dat[493] = 8'b00000000;
dat[494] = 8'b00000000;
dat[495] = 8'b00000000;
dat[496] = 8'b00000000;
dat[497] = 8'b00000000;
dat[498] = 8'b00000000;
dat[499] = 8'b00000000;
dat[500] = 8'b00000000;
dat[501] = 8'b00000000;
dat[502] = 8'b00000000;
dat[503] = 8'b00000000;
dat[504] = 8'b00000000;
dat[505] = 8'b00000000;
dat[506] = 8'b00000000;
dat[507] = 8'b00000000;
dat[508] = 8'b00000000;
dat[509] = 8'b00000000;
dat[510] = 8'b00000000;
dat[511] = 8'b00000000;
dat[512] = 8'b00000000;
dat[513] = 8'b00000000;
dat[514] = 8'b00000000;
dat[515] = 8'b00000000;
dat[516] = 8'b00000000;
dat[517] = 8'b00000000;
dat[518] = 8'b00000000;
dat[519] = 8'b00000000;
dat[520] = 8'b00000000;
dat[521] = 8'b00000000;
dat[522] = 8'b00000000;
dat[523] = 8'b00000000;
dat[524] = 8'b00000000;
dat[525] = 8'b00000000;
dat[526] = 8'b00000000;
dat[527] = 8'b00000000;
dat[528] = 8'b00000000;
dat[529] = 8'b00000000;
dat[530] = 8'b00000000;
dat[531] = 8'b00000000;
dat[532] = 8'b00000000;
dat[533] = 8'b00000000;
dat[534] = 8'b00000000;
dat[535] = 8'b00000000;
dat[536] = 8'b00000000;
dat[537] = 8'b00000000;
dat[538] = 8'b00000000;
dat[539] = 8'b00000000;
dat[540] = 8'b00000000;
dat[541] = 8'b00000000;
dat[542] = 8'b00000000;
dat[543] = 8'b00000000;
dat[544] = 8'b00000000;
dat[545] = 8'b00000000;
dat[546] = 8'b00000000;
dat[547] = 8'b00000000;
dat[548] = 8'b00000000;
dat[549] = 8'b00000000;
dat[550] = 8'b00000000;
dat[551] = 8'b00000000;
dat[552] = 8'b00000000;
dat[553] = 8'b00000000;
dat[554] = 8'b00000000;
dat[555] = 8'b00000000;
dat[556] = 8'b00000000;
dat[557] = 8'b00000000;
dat[558] = 8'b00000000;
dat[559] = 8'b00000000;
dat[560] = 8'b00000000;
dat[561] = 8'b00000000;
dat[562] = 8'b00000000;
dat[563] = 8'b00000000;
dat[564] = 8'b00000000;
dat[565] = 8'b00000000;
dat[566] = 8'b00000000;
dat[567] = 8'b00000000;
dat[568] = 8'b00000000;
dat[569] = 8'b00000000;
dat[570] = 8'b00000000;
dat[571] = 8'b00000000;
dat[572] = 8'b00000000;
dat[573] = 8'b00000000;
dat[574] = 8'b00000000;
dat[575] = 8'b00000000;
dat[576] = 8'b00000000;
dat[577] = 8'b00000000;
dat[578] = 8'b00000000;
dat[579] = 8'b00000000;
dat[580] = 8'b00000000;
dat[581] = 8'b00000000;
dat[582] = 8'b00000000;
dat[583] = 8'b00000000;
dat[584] = 8'b00000000;
dat[585] = 8'b00000000;
dat[586] = 8'b00000000;
dat[587] = 8'b00000000;
dat[588] = 8'b00000000;
dat[589] = 8'b00000000;
dat[590] = 8'b00000000;
dat[591] = 8'b00000000;
dat[592] = 8'b00000000;
dat[593] = 8'b00000000;
dat[594] = 8'b00000000;
dat[595] = 8'b00000000;
dat[596] = 8'b00000000;
dat[597] = 8'b00000000;
dat[598] = 8'b00000000;
dat[599] = 8'b00000000;
dat[600] = 8'b00000000;
dat[601] = 8'b00000000;
dat[602] = 8'b00000000;
dat[603] = 8'b00000000;
dat[604] = 8'b00000000;
dat[605] = 8'b00000000;
dat[606] = 8'b00000000;
dat[607] = 8'b00000000;
dat[608] = 8'b00000000;
dat[609] = 8'b00000000;
dat[610] = 8'b00000000;
dat[611] = 8'b00000000;
dat[612] = 8'b00000000;
dat[613] = 8'b00000000;
dat[614] = 8'b00000000;
dat[615] = 8'b00000000;
dat[616] = 8'b00000000;
dat[617] = 8'b00000000;
dat[618] = 8'b00000000;
dat[619] = 8'b00000000;
dat[620] = 8'b00000000;
dat[621] = 8'b00000000;
dat[622] = 8'b00000000;
dat[623] = 8'b00000000;
dat[624] = 8'b00000000;
dat[625] = 8'b00000000;
dat[626] = 8'b00000000;
dat[627] = 8'b00000000;
dat[628] = 8'b00000000;
dat[629] = 8'b00000000;
dat[630] = 8'b00000000;
dat[631] = 8'b00000000;
dat[632] = 8'b00000000;
dat[633] = 8'b00000000;
dat[634] = 8'b00000000;
dat[635] = 8'b00000000;
dat[636] = 8'b00000000;
dat[637] = 8'b00000000;
dat[638] = 8'b00000000;
dat[639] = 8'b00000000;
dat[640] = 8'b00000000;
dat[641] = 8'b00000000;
dat[642] = 8'b00000000;
dat[643] = 8'b00000000;
dat[644] = 8'b00000000;
dat[645] = 8'b00000000;
dat[646] = 8'b00000000;
dat[647] = 8'b00000000;
dat[648] = 8'b00000000;
dat[649] = 8'b00000000;
dat[650] = 8'b00000000;
dat[651] = 8'b00000000;
dat[652] = 8'b00000000;
dat[653] = 8'b00000000;
dat[654] = 8'b00000000;
dat[655] = 8'b00000000;
dat[656] = 8'b00000000;
dat[657] = 8'b00000000;
dat[658] = 8'b00000000;
dat[659] = 8'b00000000;
dat[660] = 8'b00000000;
dat[661] = 8'b00000000;
dat[662] = 8'b00000000;
dat[663] = 8'b00000000;
dat[664] = 8'b00000000;
dat[665] = 8'b00000000;
dat[666] = 8'b00000000;
dat[667] = 8'b00000000;
dat[668] = 8'b00000000;
dat[669] = 8'b00000000;
dat[670] = 8'b00000000;
dat[671] = 8'b00000000;
dat[672] = 8'b00000000;
dat[673] = 8'b00000000;
dat[674] = 8'b00000000;
dat[675] = 8'b00000000;
dat[676] = 8'b00000000;
dat[677] = 8'b00000000;
dat[678] = 8'b00000000;
dat[679] = 8'b00000000;
dat[680] = 8'b00000000;
dat[681] = 8'b00000000;
dat[682] = 8'b00000000;
dat[683] = 8'b00000000;
dat[684] = 8'b00000000;
dat[685] = 8'b00000000;
dat[686] = 8'b00000000;
dat[687] = 8'b00000000;
dat[688] = 8'b00000000;
dat[689] = 8'b00000000;
dat[690] = 8'b00000000;
dat[691] = 8'b00000000;
dat[692] = 8'b00000000;
dat[693] = 8'b00000000;
dat[694] = 8'b00000000;
dat[695] = 8'b00000000;
dat[696] = 8'b00000000;
dat[697] = 8'b00000000;
dat[698] = 8'b00000000;
dat[699] = 8'b00000000;
dat[700] = 8'b00000000;
dat[701] = 8'b00000000;
dat[702] = 8'b00000000;
dat[703] = 8'b00000000;
dat[704] = 8'b00000000;
dat[705] = 8'b00000000;
dat[706] = 8'b00000000;
dat[707] = 8'b00000000;
dat[708] = 8'b00000000;
dat[709] = 8'b00000000;
dat[710] = 8'b00000000;
dat[711] = 8'b00000000;
dat[712] = 8'b00000000;
dat[713] = 8'b00000000;
dat[714] = 8'b00000000;
dat[715] = 8'b00000000;
dat[716] = 8'b00000000;
dat[717] = 8'b00000000;
dat[718] = 8'b00000000;
dat[719] = 8'b00000000;
dat[720] = 8'b00000000;
dat[721] = 8'b00000000;
dat[722] = 8'b00000000;
dat[723] = 8'b00000000;
dat[724] = 8'b00000000;
dat[725] = 8'b00000000;
dat[726] = 8'b00000000;
dat[727] = 8'b00000000;
dat[728] = 8'b00000000;
dat[729] = 8'b00000000;
dat[730] = 8'b00000000;
dat[731] = 8'b00000000;
dat[732] = 8'b00000000;
dat[733] = 8'b00000000;
dat[734] = 8'b00000000;
dat[735] = 8'b00000000;
dat[736] = 8'b00000000;
dat[737] = 8'b00000000;
dat[738] = 8'b00000000;
dat[739] = 8'b00000000;
dat[740] = 8'b00000000;
dat[741] = 8'b00000000;
dat[742] = 8'b00000000;
dat[743] = 8'b00000000;
dat[744] = 8'b00000000;
dat[745] = 8'b00000000;
dat[746] = 8'b00000000;
dat[747] = 8'b00000000;
dat[748] = 8'b00000000;
dat[749] = 8'b00000000;
dat[750] = 8'b00000000;
dat[751] = 8'b00000000;
dat[752] = 8'b00000000;
dat[753] = 8'b00000000;
dat[754] = 8'b00000000;
dat[755] = 8'b00000000;
dat[756] = 8'b00000000;
dat[757] = 8'b00000000;
dat[758] = 8'b00000000;
dat[759] = 8'b00000000;
dat[760] = 8'b00000000;
dat[761] = 8'b00000000;
dat[762] = 8'b00000000;
dat[763] = 8'b00000000;
dat[764] = 8'b00000000;
dat[765] = 8'b00000000;
dat[766] = 8'b00000000;
dat[767] = 8'b00000000;
dat[768] = 8'b00000000;
dat[769] = 8'b00000000;
dat[770] = 8'b00000000;
dat[771] = 8'b00000000;
dat[772] = 8'b00000000;
dat[773] = 8'b00000000;
dat[774] = 8'b00000000;
dat[775] = 8'b00000000;
dat[776] = 8'b00000000;
dat[777] = 8'b00000000;
dat[778] = 8'b00000000;
dat[779] = 8'b00000000;
dat[780] = 8'b00000000;
dat[781] = 8'b00000000;
dat[782] = 8'b00000000;
dat[783] = 8'b00000000;
dat[784] = 8'b00000000;
dat[785] = 8'b00000000;
dat[786] = 8'b00000000;
dat[787] = 8'b00000000;
dat[788] = 8'b00000000;
dat[789] = 8'b00000000;
dat[790] = 8'b00000000;
dat[791] = 8'b00000000;
dat[792] = 8'b00000000;
dat[793] = 8'b00000000;
dat[794] = 8'b00000000;
dat[795] = 8'b00000000;
dat[796] = 8'b00000000;
dat[797] = 8'b00000000;
dat[798] = 8'b00000000;
dat[799] = 8'b00000000;
dat[800] = 8'b00000000;
dat[801] = 8'b00000000;
dat[802] = 8'b00000000;
dat[803] = 8'b00000000;
dat[804] = 8'b00000000;
dat[805] = 8'b00000000;
dat[806] = 8'b00000000;
dat[807] = 8'b00000000;
dat[808] = 8'b00000000;
dat[809] = 8'b00000000;
dat[810] = 8'b00000000;
dat[811] = 8'b00000000;
dat[812] = 8'b00000000;
dat[813] = 8'b00000000;
dat[814] = 8'b00000000;
dat[815] = 8'b00000000;
dat[816] = 8'b00000000;
dat[817] = 8'b00000000;
dat[818] = 8'b00000000;
dat[819] = 8'b00000000;
dat[820] = 8'b00000000;
dat[821] = 8'b00000000;
dat[822] = 8'b00000000;
dat[823] = 8'b00000000;
dat[824] = 8'b00000000;
dat[825] = 8'b00000000;
dat[826] = 8'b00000000;
dat[827] = 8'b00000000;
dat[828] = 8'b00000000;
dat[829] = 8'b00000000;
dat[830] = 8'b00000000;
dat[831] = 8'b00000000;
dat[832] = 8'b00000000;
dat[833] = 8'b00000000;
dat[834] = 8'b00000000;
dat[835] = 8'b00000000;
dat[836] = 8'b00000000;
dat[837] = 8'b00000000;
dat[838] = 8'b00000000;
dat[839] = 8'b00000000;
dat[840] = 8'b00000000;
dat[841] = 8'b00000000;
dat[842] = 8'b00000000;
dat[843] = 8'b00000000;
dat[844] = 8'b00000000;
dat[845] = 8'b00000000;
dat[846] = 8'b00000000;
dat[847] = 8'b00000000;
dat[848] = 8'b00000000;
dat[849] = 8'b00000000;
dat[850] = 8'b00000000;
dat[851] = 8'b00000000;
dat[852] = 8'b00000000;
dat[853] = 8'b00000000;
dat[854] = 8'b00000000;
dat[855] = 8'b00000000;
dat[856] = 8'b00000000;
dat[857] = 8'b00000000;
dat[858] = 8'b00000000;
dat[859] = 8'b00000000;
dat[860] = 8'b00000000;
dat[861] = 8'b00000000;
dat[862] = 8'b00000000;
dat[863] = 8'b00000000;
dat[864] = 8'b00000000;
dat[865] = 8'b00000000;
dat[866] = 8'b00000000;
dat[867] = 8'b00000000;
dat[868] = 8'b00000000;
dat[869] = 8'b00000000;
dat[870] = 8'b00000000;
dat[871] = 8'b00000000;
dat[872] = 8'b00000000;
dat[873] = 8'b00000000;
dat[874] = 8'b00000000;
dat[875] = 8'b00000000;
dat[876] = 8'b00000000;
dat[877] = 8'b00000000;
dat[878] = 8'b00000000;
dat[879] = 8'b00000000;
dat[880] = 8'b00000000;
dat[881] = 8'b00000000;
dat[882] = 8'b00000000;
dat[883] = 8'b00000000;
dat[884] = 8'b00000000;
dat[885] = 8'b00000000;
dat[886] = 8'b00000000;
dat[887] = 8'b00000000;
dat[888] = 8'b00000000;
dat[889] = 8'b00000000;
dat[890] = 8'b00000000;
dat[891] = 8'b00000000;
dat[892] = 8'b00000000;
dat[893] = 8'b00000000;
dat[894] = 8'b00000000;
dat[895] = 8'b00000000;
dat[896] = 8'b00000000;
dat[897] = 8'b00000000;
dat[898] = 8'b00000000;
dat[899] = 8'b00000000;
dat[900] = 8'b00000000;
dat[901] = 8'b00000000;
dat[902] = 8'b00000000;
dat[903] = 8'b00000000;
dat[904] = 8'b00000000;
dat[905] = 8'b00000000;
dat[906] = 8'b00000000;
dat[907] = 8'b00000000;
dat[908] = 8'b00000000;
dat[909] = 8'b00000000;
dat[910] = 8'b00000000;
dat[911] = 8'b00000000;
dat[912] = 8'b00000000;
dat[913] = 8'b00000000;
dat[914] = 8'b00000000;
dat[915] = 8'b00000000;
dat[916] = 8'b00000000;
dat[917] = 8'b00000000;
dat[918] = 8'b00000000;
dat[919] = 8'b00000000;
dat[920] = 8'b00000000;
dat[921] = 8'b00000000;
dat[922] = 8'b00000000;
dat[923] = 8'b00000000;
dat[924] = 8'b00000000;
dat[925] = 8'b00000000;
dat[926] = 8'b00000000;
dat[927] = 8'b00000000;
dat[928] = 8'b00000000;
dat[929] = 8'b00000000;
dat[930] = 8'b00000000;
dat[931] = 8'b00000000;
dat[932] = 8'b00000000;
dat[933] = 8'b00000000;
dat[934] = 8'b00000000;
dat[935] = 8'b00000000;
dat[936] = 8'b00000000;
dat[937] = 8'b00000000;
dat[938] = 8'b00000000;
dat[939] = 8'b00000000;
dat[940] = 8'b00000000;
dat[941] = 8'b00000000;
dat[942] = 8'b00000000;
dat[943] = 8'b00000000;
dat[944] = 8'b00000000;
dat[945] = 8'b00000000;
dat[946] = 8'b00000000;
dat[947] = 8'b00000000;
dat[948] = 8'b00000000;
dat[949] = 8'b00000000;
dat[950] = 8'b00000000;
dat[951] = 8'b00000000;
dat[952] = 8'b00000000;
dat[953] = 8'b00000000;
dat[954] = 8'b00000000;
dat[955] = 8'b00000000;
dat[956] = 8'b00000000;
dat[957] = 8'b00000000;
dat[958] = 8'b00000000;
dat[959] = 8'b00000000;
dat[960] = 8'b00000000;
dat[961] = 8'b00000000;
dat[962] = 8'b00000000;
dat[963] = 8'b00000000;
dat[964] = 8'b00000000;
dat[965] = 8'b00000000;
dat[966] = 8'b00000000;
dat[967] = 8'b00000000;
dat[968] = 8'b00000000;
dat[969] = 8'b00000000;
dat[970] = 8'b00000000;
dat[971] = 8'b00000000;
dat[972] = 8'b00000000;
dat[973] = 8'b00000000;
dat[974] = 8'b00000000;
dat[975] = 8'b00000000;
dat[976] = 8'b00000000;
dat[977] = 8'b00000000;
dat[978] = 8'b00000000;
dat[979] = 8'b00000000;
dat[980] = 8'b00000000;
dat[981] = 8'b00000000;
dat[982] = 8'b00000000;
dat[983] = 8'b00000000;
dat[984] = 8'b00000000;
dat[985] = 8'b00000000;
dat[986] = 8'b00000000;
dat[987] = 8'b00000000;
dat[988] = 8'b00000000;
dat[989] = 8'b00000000;
dat[990] = 8'b00000000;
dat[991] = 8'b00000000;
dat[992] = 8'b00000000;
dat[993] = 8'b00000000;
dat[994] = 8'b00000000;
dat[995] = 8'b00000000;
dat[996] = 8'b00000000;
dat[997] = 8'b00000000;
dat[998] = 8'b00000000;
dat[999] = 8'b00000000;
dat[1000] = 8'b00000000;
dat[1001] = 8'b00000000;
dat[1002] = 8'b00000000;
dat[1003] = 8'b00000000;
dat[1004] = 8'b00000000;
dat[1005] = 8'b00000000;
dat[1006] = 8'b00000000;
dat[1007] = 8'b00000000;
dat[1008] = 8'b00000000;
dat[1009] = 8'b00000000;
dat[1010] = 8'b00000000;
dat[1011] = 8'b00000000;
dat[1012] = 8'b00000000;
dat[1013] = 8'b00000000;
dat[1014] = 8'b00000000;
dat[1015] = 8'b00000000;
dat[1016] = 8'b00000000;
dat[1017] = 8'b00000000;
dat[1018] = 8'b00000000;
dat[1019] = 8'b00000000;
dat[1020] = 8'b00000000;
dat[1021] = 8'b00000000;
dat[1022] = 8'b00000000;
dat[1023] = 8'b00000000;
dat[1024] = 8'b00000000;
dat[1025] = 8'b00000000;
dat[1026] = 8'b00000000;
dat[1027] = 8'b00000000;
dat[1028] = 8'b00000000;
dat[1029] = 8'b00000000;
dat[1030] = 8'b00000000;
dat[1031] = 8'b00000000;
dat[1032] = 8'b00000000;
dat[1033] = 8'b00000000;
dat[1034] = 8'b00000000;
dat[1035] = 8'b00000000;
dat[1036] = 8'b00000000;
dat[1037] = 8'b00000000;
dat[1038] = 8'b00000000;
dat[1039] = 8'b00000000;
dat[1040] = 8'b00000000;
dat[1041] = 8'b00000000;
dat[1042] = 8'b00000000;
dat[1043] = 8'b00000000;
dat[1044] = 8'b00000000;
dat[1045] = 8'b00000000;
dat[1046] = 8'b00000000;
dat[1047] = 8'b00000000;
dat[1048] = 8'b00000000;
dat[1049] = 8'b00000000;
dat[1050] = 8'b00000000;
dat[1051] = 8'b00000000;
dat[1052] = 8'b00000000;
dat[1053] = 8'b00000000;
dat[1054] = 8'b00000000;
dat[1055] = 8'b00000000;
dat[1056] = 8'b00000000;
dat[1057] = 8'b00000000;
dat[1058] = 8'b00000000;
dat[1059] = 8'b00000000;
dat[1060] = 8'b00000000;
dat[1061] = 8'b00000000;
dat[1062] = 8'b00000000;
dat[1063] = 8'b00000000;
dat[1064] = 8'b00000000;
dat[1065] = 8'b00000000;
dat[1066] = 8'b00000000;
dat[1067] = 8'b00000000;
dat[1068] = 8'b00000000;
dat[1069] = 8'b00000000;
dat[1070] = 8'b00000000;
dat[1071] = 8'b00000000;
dat[1072] = 8'b00000000;
dat[1073] = 8'b00000000;
dat[1074] = 8'b00000000;
dat[1075] = 8'b00000000;
dat[1076] = 8'b00000000;
dat[1077] = 8'b00000000;
dat[1078] = 8'b00000000;
dat[1079] = 8'b00000000;
dat[1080] = 8'b00000000;
dat[1081] = 8'b00000000;
dat[1082] = 8'b00000000;
dat[1083] = 8'b00000000;
dat[1084] = 8'b00000000;
dat[1085] = 8'b00000000;
dat[1086] = 8'b00000000;
dat[1087] = 8'b00000000;
dat[1088] = 8'b00000000;
dat[1089] = 8'b00000000;
dat[1090] = 8'b00000000;
dat[1091] = 8'b00000000;
dat[1092] = 8'b00000000;
dat[1093] = 8'b00000000;
dat[1094] = 8'b00000000;
dat[1095] = 8'b00000000;
dat[1096] = 8'b00000000;
dat[1097] = 8'b00000000;
dat[1098] = 8'b00000000;
dat[1099] = 8'b00000000;
dat[1100] = 8'b00000000;
dat[1101] = 8'b00000000;
dat[1102] = 8'b00000000;
dat[1103] = 8'b00000000;
dat[1104] = 8'b00000000;
dat[1105] = 8'b00000000;
dat[1106] = 8'b00000000;
dat[1107] = 8'b00000000;
dat[1108] = 8'b00000000;
dat[1109] = 8'b00000000;
dat[1110] = 8'b00000000;
dat[1111] = 8'b00000000;
dat[1112] = 8'b00000000;
dat[1113] = 8'b00000000;
dat[1114] = 8'b00000000;
dat[1115] = 8'b00000000;
dat[1116] = 8'b00000000;
dat[1117] = 8'b00000000;
dat[1118] = 8'b00000000;
dat[1119] = 8'b00000000;
dat[1120] = 8'b00000000;
dat[1121] = 8'b00000000;
dat[1122] = 8'b00000000;
dat[1123] = 8'b00000000;
dat[1124] = 8'b00000000;
dat[1125] = 8'b00000000;
dat[1126] = 8'b00000000;
dat[1127] = 8'b00000000;
dat[1128] = 8'b00000000;
dat[1129] = 8'b00000000;
dat[1130] = 8'b00000000;
dat[1131] = 8'b00000000;
dat[1132] = 8'b00000000;
dat[1133] = 8'b00000000;
dat[1134] = 8'b00000000;
dat[1135] = 8'b00000000;
dat[1136] = 8'b00000000;
dat[1137] = 8'b00000000;
dat[1138] = 8'b00000000;
dat[1139] = 8'b00000000;
dat[1140] = 8'b00000000;
dat[1141] = 8'b00000000;
dat[1142] = 8'b00000000;
dat[1143] = 8'b00000000;
dat[1144] = 8'b00000000;
dat[1145] = 8'b00000000;
dat[1146] = 8'b00000000;
dat[1147] = 8'b00000000;
dat[1148] = 8'b00000000;
dat[1149] = 8'b00000000;
dat[1150] = 8'b00000000;
dat[1151] = 8'b00000000;
dat[1152] = 8'b00000000;
dat[1153] = 8'b00000000;
dat[1154] = 8'b00000000;
dat[1155] = 8'b00000000;
dat[1156] = 8'b00000000;
dat[1157] = 8'b00000000;
dat[1158] = 8'b00000000;
dat[1159] = 8'b00000000;
dat[1160] = 8'b00000000;
dat[1161] = 8'b00000000;
dat[1162] = 8'b00000000;
dat[1163] = 8'b00000000;
dat[1164] = 8'b00000000;
dat[1165] = 8'b00000000;
dat[1166] = 8'b00000000;
dat[1167] = 8'b00000000;
dat[1168] = 8'b00000000;
dat[1169] = 8'b00000000;
dat[1170] = 8'b00000000;
dat[1171] = 8'b00000000;
dat[1172] = 8'b00000000;
dat[1173] = 8'b00000000;
dat[1174] = 8'b00000000;
dat[1175] = 8'b00000000;
dat[1176] = 8'b00000000;
dat[1177] = 8'b00000000;
dat[1178] = 8'b00000000;
dat[1179] = 8'b00000000;
dat[1180] = 8'b00000000;
dat[1181] = 8'b00000000;
dat[1182] = 8'b00000000;
dat[1183] = 8'b00000000;
dat[1184] = 8'b00000000;
dat[1185] = 8'b00000000;
dat[1186] = 8'b00000000;
dat[1187] = 8'b00000000;
dat[1188] = 8'b00000000;
dat[1189] = 8'b00000000;
dat[1190] = 8'b00000000;
dat[1191] = 8'b00000000;
dat[1192] = 8'b00000000;
dat[1193] = 8'b00000000;
dat[1194] = 8'b00000000;
dat[1195] = 8'b00000000;
dat[1196] = 8'b00000000;
dat[1197] = 8'b00000000;
dat[1198] = 8'b00000000;
dat[1199] = 8'b00000000;
dat[1200] = 8'b00000000;
dat[1201] = 8'b00000000;
dat[1202] = 8'b00000000;
dat[1203] = 8'b00000000;
dat[1204] = 8'b00000000;
dat[1205] = 8'b00000000;
dat[1206] = 8'b00000000;
dat[1207] = 8'b00000000;
dat[1208] = 8'b00000000;
dat[1209] = 8'b00000000;
dat[1210] = 8'b00000000;
dat[1211] = 8'b00000000;
dat[1212] = 8'b00000000;
dat[1213] = 8'b00000000;
dat[1214] = 8'b00000000;
dat[1215] = 8'b00000000;
dat[1216] = 8'b00000000;
dat[1217] = 8'b00000000;
dat[1218] = 8'b00000000;
dat[1219] = 8'b00000000;
dat[1220] = 8'b00000000;
dat[1221] = 8'b00000000;
dat[1222] = 8'b00000000;
dat[1223] = 8'b00000000;
dat[1224] = 8'b00000000;
dat[1225] = 8'b00000000;
dat[1226] = 8'b00000000;
dat[1227] = 8'b00000000;
dat[1228] = 8'b00000000;
dat[1229] = 8'b00000000;
dat[1230] = 8'b00000000;
dat[1231] = 8'b00000000;
dat[1232] = 8'b00000000;
dat[1233] = 8'b00000000;
dat[1234] = 8'b00000000;
dat[1235] = 8'b00000000;
dat[1236] = 8'b00000000;
dat[1237] = 8'b00000000;
dat[1238] = 8'b00000000;
dat[1239] = 8'b00000000;
dat[1240] = 8'b00000000;
dat[1241] = 8'b00000000;
dat[1242] = 8'b00000000;
dat[1243] = 8'b00000000;
dat[1244] = 8'b00000000;
dat[1245] = 8'b00000000;
dat[1246] = 8'b00000000;
dat[1247] = 8'b00000000;
dat[1248] = 8'b00000000;
dat[1249] = 8'b00000000;
dat[1250] = 8'b00000000;
dat[1251] = 8'b00000000;
dat[1252] = 8'b00000000;
dat[1253] = 8'b00000000;
dat[1254] = 8'b00000000;
dat[1255] = 8'b00000000;
dat[1256] = 8'b00000000;
dat[1257] = 8'b00000000;
dat[1258] = 8'b00000000;
dat[1259] = 8'b00000000;
dat[1260] = 8'b00000000;
dat[1261] = 8'b00000000;
dat[1262] = 8'b00000000;
dat[1263] = 8'b00000000;
dat[1264] = 8'b00000000;
dat[1265] = 8'b00000000;
dat[1266] = 8'b00000000;
dat[1267] = 8'b00000000;
dat[1268] = 8'b00000000;
dat[1269] = 8'b00000000;
dat[1270] = 8'b00000000;
dat[1271] = 8'b00000000;
dat[1272] = 8'b00000000;
dat[1273] = 8'b00000000;
dat[1274] = 8'b00000000;
dat[1275] = 8'b00000000;
dat[1276] = 8'b00000000;
dat[1277] = 8'b00000000;
dat[1278] = 8'b00000000;
dat[1279] = 8'b00000000;
dat[1280] = 8'b00000000;
dat[1281] = 8'b00000000;
dat[1282] = 8'b00000000;
dat[1283] = 8'b00000000;
dat[1284] = 8'b00000000;
dat[1285] = 8'b00000000;
dat[1286] = 8'b00000000;
dat[1287] = 8'b00000000;
dat[1288] = 8'b00000000;
dat[1289] = 8'b00000000;
dat[1290] = 8'b00000000;
dat[1291] = 8'b00000000;
dat[1292] = 8'b00000000;
dat[1293] = 8'b00000000;
dat[1294] = 8'b00000000;
dat[1295] = 8'b00000000;
dat[1296] = 8'b00000000;
dat[1297] = 8'b00000000;
dat[1298] = 8'b00000000;
dat[1299] = 8'b00000000;
dat[1300] = 8'b00000000;
dat[1301] = 8'b00000000;
dat[1302] = 8'b00000000;
dat[1303] = 8'b00000000;
dat[1304] = 8'b00000000;
dat[1305] = 8'b00000000;
dat[1306] = 8'b00000000;
dat[1307] = 8'b00000000;
dat[1308] = 8'b00000000;
dat[1309] = 8'b00000000;
dat[1310] = 8'b00000000;
dat[1311] = 8'b00000000;
dat[1312] = 8'b00000000;
dat[1313] = 8'b00000000;
dat[1314] = 8'b00000000;
dat[1315] = 8'b00000000;
dat[1316] = 8'b00000000;
dat[1317] = 8'b00000000;
dat[1318] = 8'b00000000;
dat[1319] = 8'b00000000;
dat[1320] = 8'b00000000;
dat[1321] = 8'b00000000;
dat[1322] = 8'b00000000;
dat[1323] = 8'b00000000;
dat[1324] = 8'b00000000;
dat[1325] = 8'b00000000;
dat[1326] = 8'b00000000;
dat[1327] = 8'b00000000;
dat[1328] = 8'b00000000;
dat[1329] = 8'b00000000;
dat[1330] = 8'b00000000;
dat[1331] = 8'b00000000;
dat[1332] = 8'b00000000;
dat[1333] = 8'b00000000;
dat[1334] = 8'b00000000;
dat[1335] = 8'b00000000;
dat[1336] = 8'b00000000;
dat[1337] = 8'b00000000;
dat[1338] = 8'b00000000;
dat[1339] = 8'b00000000;
dat[1340] = 8'b00000000;
dat[1341] = 8'b00000000;
dat[1342] = 8'b00000000;
dat[1343] = 8'b00000000;
dat[1344] = 8'b00000000;
dat[1345] = 8'b00000000;
dat[1346] = 8'b00000000;
dat[1347] = 8'b00000000;
dat[1348] = 8'b00000000;
dat[1349] = 8'b00000000;
dat[1350] = 8'b00000000;
dat[1351] = 8'b00000000;
dat[1352] = 8'b00000000;
dat[1353] = 8'b00000000;
dat[1354] = 8'b00000000;
dat[1355] = 8'b00000000;
dat[1356] = 8'b00000000;
dat[1357] = 8'b00000000;
dat[1358] = 8'b00000000;
dat[1359] = 8'b00000000;
dat[1360] = 8'b00000000;
dat[1361] = 8'b00000000;
dat[1362] = 8'b00000000;
dat[1363] = 8'b00000000;
dat[1364] = 8'b00000000;
dat[1365] = 8'b00000000;
dat[1366] = 8'b00000000;
dat[1367] = 8'b00000000;
dat[1368] = 8'b00000000;
dat[1369] = 8'b00000000;
dat[1370] = 8'b00000000;
dat[1371] = 8'b00000000;
dat[1372] = 8'b00000000;
dat[1373] = 8'b00000000;
dat[1374] = 8'b00000000;
dat[1375] = 8'b00000000;
dat[1376] = 8'b00000000;
dat[1377] = 8'b00000000;
dat[1378] = 8'b00000000;
dat[1379] = 8'b00000000;
dat[1380] = 8'b00000000;
dat[1381] = 8'b00000000;
dat[1382] = 8'b00000000;
dat[1383] = 8'b00000000;
dat[1384] = 8'b00000000;
dat[1385] = 8'b00000000;
dat[1386] = 8'b00000000;
dat[1387] = 8'b00000000;
dat[1388] = 8'b00000000;
dat[1389] = 8'b00000000;
dat[1390] = 8'b00000000;
dat[1391] = 8'b00000000;
dat[1392] = 8'b00000000;
dat[1393] = 8'b00000000;
dat[1394] = 8'b00000000;
dat[1395] = 8'b00000000;
dat[1396] = 8'b00000000;
dat[1397] = 8'b00000000;
dat[1398] = 8'b00000000;
dat[1399] = 8'b00000000;
dat[1400] = 8'b00000000;
dat[1401] = 8'b00000000;
dat[1402] = 8'b00000000;
dat[1403] = 8'b00000000;
dat[1404] = 8'b00000000;
dat[1405] = 8'b00000000;
dat[1406] = 8'b00000000;
dat[1407] = 8'b00000000;
dat[1408] = 8'b00000000;
dat[1409] = 8'b00000000;
dat[1410] = 8'b00000000;
dat[1411] = 8'b00000000;
dat[1412] = 8'b00000000;
dat[1413] = 8'b00000000;
dat[1414] = 8'b00000000;
dat[1415] = 8'b00000000;
dat[1416] = 8'b00000000;
dat[1417] = 8'b00000000;
dat[1418] = 8'b00000000;
dat[1419] = 8'b00000000;
dat[1420] = 8'b00000000;
dat[1421] = 8'b00000000;
dat[1422] = 8'b00000000;
dat[1423] = 8'b00000000;
dat[1424] = 8'b00000000;
dat[1425] = 8'b00000000;
dat[1426] = 8'b00000000;
dat[1427] = 8'b00000000;
dat[1428] = 8'b00000000;
dat[1429] = 8'b00000000;
dat[1430] = 8'b00000000;
dat[1431] = 8'b00000000;
dat[1432] = 8'b00000000;
dat[1433] = 8'b00000000;
dat[1434] = 8'b00000000;
dat[1435] = 8'b00000000;
dat[1436] = 8'b00000000;
dat[1437] = 8'b00000000;
dat[1438] = 8'b00000000;
dat[1439] = 8'b00000000;
dat[1440] = 8'b00000000;
dat[1441] = 8'b00000000;
dat[1442] = 8'b00000000;
dat[1443] = 8'b00000000;
dat[1444] = 8'b00000000;
dat[1445] = 8'b00000000;
dat[1446] = 8'b00000000;
dat[1447] = 8'b00000000;
dat[1448] = 8'b00000000;
dat[1449] = 8'b00000000;
dat[1450] = 8'b00000000;
dat[1451] = 8'b00000000;
dat[1452] = 8'b00000000;
dat[1453] = 8'b00000000;
dat[1454] = 8'b00000000;
dat[1455] = 8'b00000000;
dat[1456] = 8'b00000000;
dat[1457] = 8'b00000000;
dat[1458] = 8'b00000000;
dat[1459] = 8'b00000000;
dat[1460] = 8'b00000000;
dat[1461] = 8'b00000000;
dat[1462] = 8'b00000000;
dat[1463] = 8'b00000000;
dat[1464] = 8'b00000000;
dat[1465] = 8'b00000000;
dat[1466] = 8'b00000000;
dat[1467] = 8'b00000000;
dat[1468] = 8'b00000000;
dat[1469] = 8'b00000000;
dat[1470] = 8'b00000000;
dat[1471] = 8'b00000000;
dat[1472] = 8'b00000000;
dat[1473] = 8'b00000000;
dat[1474] = 8'b00000000;
dat[1475] = 8'b00000000;
dat[1476] = 8'b00000000;
dat[1477] = 8'b00000000;
dat[1478] = 8'b00000000;
dat[1479] = 8'b00000000;
dat[1480] = 8'b00000000;
dat[1481] = 8'b00000000;
dat[1482] = 8'b00000000;
dat[1483] = 8'b00000000;
dat[1484] = 8'b00000000;
dat[1485] = 8'b00000000;
dat[1486] = 8'b00000000;
dat[1487] = 8'b00000000;
dat[1488] = 8'b00000000;
dat[1489] = 8'b00000000;
dat[1490] = 8'b00000000;
dat[1491] = 8'b00000000;
dat[1492] = 8'b00000000;
dat[1493] = 8'b00000000;
dat[1494] = 8'b00000000;
dat[1495] = 8'b00000000;
dat[1496] = 8'b00000000;
dat[1497] = 8'b00000000;
dat[1498] = 8'b00000000;
dat[1499] = 8'b00000000;
dat[1500] = 8'b00000000;
dat[1501] = 8'b00000000;
dat[1502] = 8'b00000000;
dat[1503] = 8'b00000000;
dat[1504] = 8'b00000000;
dat[1505] = 8'b00000000;
dat[1506] = 8'b00000000;
dat[1507] = 8'b00000000;
dat[1508] = 8'b00000000;
dat[1509] = 8'b00000000;
dat[1510] = 8'b00000000;
dat[1511] = 8'b00000000;
dat[1512] = 8'b00000000;
dat[1513] = 8'b00000000;
dat[1514] = 8'b00000000;
dat[1515] = 8'b00000000;
dat[1516] = 8'b00000000;
dat[1517] = 8'b00000000;
dat[1518] = 8'b00000000;
dat[1519] = 8'b00000000;
dat[1520] = 8'b00000000;
dat[1521] = 8'b00000000;
dat[1522] = 8'b00000000;
dat[1523] = 8'b00000000;
dat[1524] = 8'b00000000;
dat[1525] = 8'b00000000;
dat[1526] = 8'b00000000;
dat[1527] = 8'b00000000;
dat[1528] = 8'b00000000;
dat[1529] = 8'b00000000;
dat[1530] = 8'b00000000;
dat[1531] = 8'b00000000;
dat[1532] = 8'b00000000;
dat[1533] = 8'b00000000;
dat[1534] = 8'b00000000;
dat[1535] = 8'b00000000;
dat[1536] = 8'b00000000;
dat[1537] = 8'b00000000;
dat[1538] = 8'b00000000;
dat[1539] = 8'b00000000;
dat[1540] = 8'b00000000;
dat[1541] = 8'b00000000;
dat[1542] = 8'b00000000;
dat[1543] = 8'b00000000;
dat[1544] = 8'b00000000;
dat[1545] = 8'b00000000;
dat[1546] = 8'b00000000;
dat[1547] = 8'b00000000;
dat[1548] = 8'b00000000;
dat[1549] = 8'b00000000;
dat[1550] = 8'b00000000;
dat[1551] = 8'b00000000;
dat[1552] = 8'b00000000;
dat[1553] = 8'b00000000;
dat[1554] = 8'b00000000;
dat[1555] = 8'b00000000;
dat[1556] = 8'b00000000;
dat[1557] = 8'b00000000;
dat[1558] = 8'b00000000;
dat[1559] = 8'b00000000;
dat[1560] = 8'b00000000;
dat[1561] = 8'b00000000;
dat[1562] = 8'b00000000;
dat[1563] = 8'b00000000;
dat[1564] = 8'b00000000;
dat[1565] = 8'b00000000;
dat[1566] = 8'b00000000;
dat[1567] = 8'b00000000;
dat[1568] = 8'b00000000;
dat[1569] = 8'b00000000;
dat[1570] = 8'b00000000;
dat[1571] = 8'b00000000;
dat[1572] = 8'b00000000;
dat[1573] = 8'b00000000;
dat[1574] = 8'b00000000;
dat[1575] = 8'b00000000;
dat[1576] = 8'b00000000;
dat[1577] = 8'b00000000;
dat[1578] = 8'b00000000;
dat[1579] = 8'b00000000;
dat[1580] = 8'b00000000;
dat[1581] = 8'b00000000;
dat[1582] = 8'b00000000;
dat[1583] = 8'b00000000;
dat[1584] = 8'b00000000;
dat[1585] = 8'b00000000;
dat[1586] = 8'b00000000;
dat[1587] = 8'b00000000;
dat[1588] = 8'b00000000;
dat[1589] = 8'b00000000;
dat[1590] = 8'b00000000;
dat[1591] = 8'b00000000;
dat[1592] = 8'b00000000;
dat[1593] = 8'b00000000;
dat[1594] = 8'b00000000;
dat[1595] = 8'b00000000;
dat[1596] = 8'b00000000;
dat[1597] = 8'b00000000;
dat[1598] = 8'b00000000;
dat[1599] = 8'b00000000;
dat[1600] = 8'b00000000;
dat[1601] = 8'b00000000;
dat[1602] = 8'b00000000;
dat[1603] = 8'b00000000;
dat[1604] = 8'b00000000;
dat[1605] = 8'b00000000;
dat[1606] = 8'b00000000;
dat[1607] = 8'b00000000;
dat[1608] = 8'b00000000;
dat[1609] = 8'b00000000;
dat[1610] = 8'b00000000;
dat[1611] = 8'b00000000;
dat[1612] = 8'b00000000;
dat[1613] = 8'b00000000;
dat[1614] = 8'b00000000;
dat[1615] = 8'b00000000;
dat[1616] = 8'b00000000;
dat[1617] = 8'b00000000;
dat[1618] = 8'b00000000;
dat[1619] = 8'b00000000;
dat[1620] = 8'b00000000;
dat[1621] = 8'b00000000;
dat[1622] = 8'b00000000;
dat[1623] = 8'b00000000;
dat[1624] = 8'b00000000;
dat[1625] = 8'b00000000;
dat[1626] = 8'b00000000;
dat[1627] = 8'b00000000;
dat[1628] = 8'b00000000;
dat[1629] = 8'b00000000;
dat[1630] = 8'b00000000;
dat[1631] = 8'b00000000;
dat[1632] = 8'b00000000;
dat[1633] = 8'b00000000;
dat[1634] = 8'b00000000;
dat[1635] = 8'b00000000;
dat[1636] = 8'b00000000;
dat[1637] = 8'b00000000;
dat[1638] = 8'b00000000;
dat[1639] = 8'b00000000;
dat[1640] = 8'b00000000;
dat[1641] = 8'b00000000;
dat[1642] = 8'b00000000;
dat[1643] = 8'b00000000;
dat[1644] = 8'b00000000;
dat[1645] = 8'b00000000;
dat[1646] = 8'b00000000;
dat[1647] = 8'b00000000;
dat[1648] = 8'b00000000;
dat[1649] = 8'b00000000;
dat[1650] = 8'b00000000;
dat[1651] = 8'b00000000;
dat[1652] = 8'b00000000;
dat[1653] = 8'b00000000;
dat[1654] = 8'b00000000;
dat[1655] = 8'b00000000;
dat[1656] = 8'b00000000;
dat[1657] = 8'b00000000;
dat[1658] = 8'b00000000;
dat[1659] = 8'b00000000;
dat[1660] = 8'b00000000;
dat[1661] = 8'b00000000;
dat[1662] = 8'b00000000;
dat[1663] = 8'b00000000;
dat[1664] = 8'b00000000;
dat[1665] = 8'b00000000;
dat[1666] = 8'b00000000;
dat[1667] = 8'b00000000;
dat[1668] = 8'b00000000;
dat[1669] = 8'b00000000;
dat[1670] = 8'b00000000;
dat[1671] = 8'b00000000;
dat[1672] = 8'b00000000;
dat[1673] = 8'b00000000;
dat[1674] = 8'b00000000;
dat[1675] = 8'b00000000;
dat[1676] = 8'b00000000;
dat[1677] = 8'b00000000;
dat[1678] = 8'b00000000;
dat[1679] = 8'b00000000;
dat[1680] = 8'b00000000;
dat[1681] = 8'b00000000;
dat[1682] = 8'b00000000;
dat[1683] = 8'b00000000;
dat[1684] = 8'b00000000;
dat[1685] = 8'b00000000;
dat[1686] = 8'b00000000;
dat[1687] = 8'b00000000;
dat[1688] = 8'b00000000;
dat[1689] = 8'b00000000;
dat[1690] = 8'b00000000;
dat[1691] = 8'b00000000;
dat[1692] = 8'b00000000;
dat[1693] = 8'b00000000;
dat[1694] = 8'b00000000;
dat[1695] = 8'b00000000;
dat[1696] = 8'b00000000;
dat[1697] = 8'b00000000;
dat[1698] = 8'b00000000;
dat[1699] = 8'b00000000;
dat[1700] = 8'b00000000;
dat[1701] = 8'b00000000;
dat[1702] = 8'b00000000;
dat[1703] = 8'b00000000;
dat[1704] = 8'b00000000;
dat[1705] = 8'b00000000;
dat[1706] = 8'b00000000;
dat[1707] = 8'b00000000;
dat[1708] = 8'b00000000;
dat[1709] = 8'b00000000;
dat[1710] = 8'b00000000;
dat[1711] = 8'b00000000;
dat[1712] = 8'b00000000;
dat[1713] = 8'b00000000;
dat[1714] = 8'b00000000;
dat[1715] = 8'b00000000;
dat[1716] = 8'b00000000;
dat[1717] = 8'b00000000;
dat[1718] = 8'b00000000;
dat[1719] = 8'b00000000;
dat[1720] = 8'b00000000;
dat[1721] = 8'b00000000;
dat[1722] = 8'b00000000;
dat[1723] = 8'b00000000;
dat[1724] = 8'b00000000;
dat[1725] = 8'b00000000;
dat[1726] = 8'b00000000;
dat[1727] = 8'b00000000;
dat[1728] = 8'b00000000;
dat[1729] = 8'b00000000;
dat[1730] = 8'b00000000;
dat[1731] = 8'b00000000;
dat[1732] = 8'b00000000;
dat[1733] = 8'b00000000;
dat[1734] = 8'b00000000;
dat[1735] = 8'b00000000;
dat[1736] = 8'b00000000;
dat[1737] = 8'b00000000;
dat[1738] = 8'b00000000;
dat[1739] = 8'b00000000;
dat[1740] = 8'b00000000;
dat[1741] = 8'b00000000;
dat[1742] = 8'b00000000;
dat[1743] = 8'b00000000;
dat[1744] = 8'b00000000;
dat[1745] = 8'b00000000;
dat[1746] = 8'b00000000;
dat[1747] = 8'b00000000;
dat[1748] = 8'b00000000;
dat[1749] = 8'b00000000;
dat[1750] = 8'b00000000;
dat[1751] = 8'b00000000;
dat[1752] = 8'b00000000;
dat[1753] = 8'b00000000;
dat[1754] = 8'b00000000;
dat[1755] = 8'b00000000;
dat[1756] = 8'b00000000;
dat[1757] = 8'b00000000;
dat[1758] = 8'b00000000;
dat[1759] = 8'b00000000;
dat[1760] = 8'b00000000;
dat[1761] = 8'b00000000;
dat[1762] = 8'b00000000;
dat[1763] = 8'b00000000;
dat[1764] = 8'b00000000;
dat[1765] = 8'b00000000;
dat[1766] = 8'b00000000;
dat[1767] = 8'b00000000;
dat[1768] = 8'b00000000;
dat[1769] = 8'b00000000;
dat[1770] = 8'b00000000;
dat[1771] = 8'b00000000;
dat[1772] = 8'b00000000;
dat[1773] = 8'b00000000;
dat[1774] = 8'b00000000;
dat[1775] = 8'b00000000;
dat[1776] = 8'b00000000;
dat[1777] = 8'b00000000;
dat[1778] = 8'b00000000;
dat[1779] = 8'b00000000;
dat[1780] = 8'b00000000;
dat[1781] = 8'b00000000;
dat[1782] = 8'b00000000;
dat[1783] = 8'b00000000;
dat[1784] = 8'b00000000;
dat[1785] = 8'b00000000;
dat[1786] = 8'b00000000;
dat[1787] = 8'b00000000;
dat[1788] = 8'b00000000;
dat[1789] = 8'b00000000;
dat[1790] = 8'b00000000;
dat[1791] = 8'b00000000;
dat[1792] = 8'b00000000;
dat[1793] = 8'b00000000;
dat[1794] = 8'b00000000;
dat[1795] = 8'b00000000;
dat[1796] = 8'b00000000;
dat[1797] = 8'b00000000;
dat[1798] = 8'b00000000;
dat[1799] = 8'b00000000;
dat[1800] = 8'b00000000;
dat[1801] = 8'b00000000;
dat[1802] = 8'b00000000;
dat[1803] = 8'b00000000;
dat[1804] = 8'b00000000;
dat[1805] = 8'b00000000;
dat[1806] = 8'b00000000;
dat[1807] = 8'b00000000;
dat[1808] = 8'b00000000;
dat[1809] = 8'b00000000;
dat[1810] = 8'b00000000;
dat[1811] = 8'b00000000;
dat[1812] = 8'b00000000;
dat[1813] = 8'b00000000;
dat[1814] = 8'b00000000;
dat[1815] = 8'b00000000;
dat[1816] = 8'b00000000;
dat[1817] = 8'b00000000;
dat[1818] = 8'b00000000;
dat[1819] = 8'b00000000;
dat[1820] = 8'b00000000;
dat[1821] = 8'b00000000;
dat[1822] = 8'b00000000;
dat[1823] = 8'b00000000;
dat[1824] = 8'b00000000;
dat[1825] = 8'b00000000;
dat[1826] = 8'b00000000;
dat[1827] = 8'b00000000;
dat[1828] = 8'b00000000;
dat[1829] = 8'b00000000;
dat[1830] = 8'b00000000;
dat[1831] = 8'b00000000;
dat[1832] = 8'b00000000;
dat[1833] = 8'b00000000;
dat[1834] = 8'b00000000;
dat[1835] = 8'b00000000;
dat[1836] = 8'b00000000;
dat[1837] = 8'b00000000;
dat[1838] = 8'b00000000;
dat[1839] = 8'b00000000;
dat[1840] = 8'b00000000;
dat[1841] = 8'b00000000;
dat[1842] = 8'b00000000;
dat[1843] = 8'b00000000;
dat[1844] = 8'b00000000;
dat[1845] = 8'b00000000;
dat[1846] = 8'b00000000;
dat[1847] = 8'b00000000;
dat[1848] = 8'b00000000;
dat[1849] = 8'b00000000;
dat[1850] = 8'b00000000;
dat[1851] = 8'b00000000;
dat[1852] = 8'b00000000;
dat[1853] = 8'b00000000;
dat[1854] = 8'b00000000;
dat[1855] = 8'b00000000;
dat[1856] = 8'b00000000;
dat[1857] = 8'b00000000;
dat[1858] = 8'b00000000;
dat[1859] = 8'b00000000;
dat[1860] = 8'b00000000;
dat[1861] = 8'b00000000;
dat[1862] = 8'b00000000;
dat[1863] = 8'b00000000;
dat[1864] = 8'b00000000;
dat[1865] = 8'b00000000;
dat[1866] = 8'b00000000;
dat[1867] = 8'b00000000;
dat[1868] = 8'b00000000;
dat[1869] = 8'b00000000;
dat[1870] = 8'b00000000;
dat[1871] = 8'b00000000;
dat[1872] = 8'b00000000;
dat[1873] = 8'b00000000;
dat[1874] = 8'b00000000;
dat[1875] = 8'b00000000;
dat[1876] = 8'b00000000;
dat[1877] = 8'b00000000;
dat[1878] = 8'b00000000;
dat[1879] = 8'b00000000;
dat[1880] = 8'b00000000;
dat[1881] = 8'b00000000;
dat[1882] = 8'b00000000;
dat[1883] = 8'b00000000;
dat[1884] = 8'b00000000;
dat[1885] = 8'b00000000;
dat[1886] = 8'b00000000;
dat[1887] = 8'b00000000;
dat[1888] = 8'b00000000;
dat[1889] = 8'b00000000;
dat[1890] = 8'b00000000;
dat[1891] = 8'b00000000;
dat[1892] = 8'b00000000;
dat[1893] = 8'b00000000;
dat[1894] = 8'b00000000;
dat[1895] = 8'b00000000;
dat[1896] = 8'b00000000;
dat[1897] = 8'b00000000;
dat[1898] = 8'b00000000;
dat[1899] = 8'b00000000;
dat[1900] = 8'b00000000;
dat[1901] = 8'b00000000;
dat[1902] = 8'b00000000;
dat[1903] = 8'b00000000;
dat[1904] = 8'b00000000;
dat[1905] = 8'b00000000;
dat[1906] = 8'b00000000;
dat[1907] = 8'b00000000;
dat[1908] = 8'b00000000;
dat[1909] = 8'b00000000;
dat[1910] = 8'b00000000;
dat[1911] = 8'b00000000;
dat[1912] = 8'b00000000;
dat[1913] = 8'b00000000;
dat[1914] = 8'b00000000;
dat[1915] = 8'b00000000;
dat[1916] = 8'b00000000;
dat[1917] = 8'b00000000;
dat[1918] = 8'b00000000;
dat[1919] = 8'b00000000;
dat[1920] = 8'b00000000;
dat[1921] = 8'b00000000;
dat[1922] = 8'b00000000;
dat[1923] = 8'b00000000;
dat[1924] = 8'b00000000;
dat[1925] = 8'b00000000;
dat[1926] = 8'b00000000;
dat[1927] = 8'b00000000;
dat[1928] = 8'b00000000;
dat[1929] = 8'b00000000;
dat[1930] = 8'b00000000;
dat[1931] = 8'b00000000;
dat[1932] = 8'b00000000;
dat[1933] = 8'b00000000;
dat[1934] = 8'b00000000;
dat[1935] = 8'b00000000;
dat[1936] = 8'b00000000;
dat[1937] = 8'b00000000;
dat[1938] = 8'b00000000;
dat[1939] = 8'b00000000;
dat[1940] = 8'b00000000;
dat[1941] = 8'b00000000;
dat[1942] = 8'b00000000;
dat[1943] = 8'b00000000;
dat[1944] = 8'b00000000;
dat[1945] = 8'b00000000;
dat[1946] = 8'b00000000;
dat[1947] = 8'b00000000;
dat[1948] = 8'b00000000;
dat[1949] = 8'b00000000;
dat[1950] = 8'b00000000;
dat[1951] = 8'b00000000;
dat[1952] = 8'b00000000;
dat[1953] = 8'b00000000;
dat[1954] = 8'b00000000;
dat[1955] = 8'b00000000;
dat[1956] = 8'b00000000;
dat[1957] = 8'b00000000;
dat[1958] = 8'b00000000;
dat[1959] = 8'b00000000;
dat[1960] = 8'b00000000;
dat[1961] = 8'b00000000;
dat[1962] = 8'b00000000;
dat[1963] = 8'b00000000;
dat[1964] = 8'b00000000;
dat[1965] = 8'b00000000;
dat[1966] = 8'b00000000;
dat[1967] = 8'b00000000;
dat[1968] = 8'b00000000;
dat[1969] = 8'b00000000;
dat[1970] = 8'b00000000;
dat[1971] = 8'b00000000;
dat[1972] = 8'b00000000;
dat[1973] = 8'b00000000;
dat[1974] = 8'b00000000;
dat[1975] = 8'b00000000;
dat[1976] = 8'b00000000;
dat[1977] = 8'b00000000;
dat[1978] = 8'b00000000;
dat[1979] = 8'b00000000;
dat[1980] = 8'b00000000;
dat[1981] = 8'b00000000;
dat[1982] = 8'b00000000;
dat[1983] = 8'b00000000;
dat[1984] = 8'b00000000;
dat[1985] = 8'b00000000;
dat[1986] = 8'b00000000;
dat[1987] = 8'b00000000;
dat[1988] = 8'b00000000;
dat[1989] = 8'b00000000;
dat[1990] = 8'b00000000;
dat[1991] = 8'b00000000;
dat[1992] = 8'b00000000;
dat[1993] = 8'b00000000;
dat[1994] = 8'b00000000;
dat[1995] = 8'b00000000;
dat[1996] = 8'b00000000;
dat[1997] = 8'b00000000;
dat[1998] = 8'b00000000;
dat[1999] = 8'b00000000;
dat[2000] = 8'b00000000;
dat[2001] = 8'b00000000;
dat[2002] = 8'b00000000;
dat[2003] = 8'b00000000;
dat[2004] = 8'b00000000;
dat[2005] = 8'b00000000;
dat[2006] = 8'b00000000;
dat[2007] = 8'b00000000;
dat[2008] = 8'b00000000;
dat[2009] = 8'b00000000;
dat[2010] = 8'b00000000;
dat[2011] = 8'b00000000;
dat[2012] = 8'b00000000;
dat[2013] = 8'b00000000;
dat[2014] = 8'b00000000;
dat[2015] = 8'b00000000;
dat[2016] = 8'b00000000;
dat[2017] = 8'b00000000;
dat[2018] = 8'b00000000;
dat[2019] = 8'b00000000;
dat[2020] = 8'b00000000;
dat[2021] = 8'b00000000;
dat[2022] = 8'b00000000;
dat[2023] = 8'b00000000;
dat[2024] = 8'b00000000;
dat[2025] = 8'b00000000;
dat[2026] = 8'b00000000;
dat[2027] = 8'b00000000;
dat[2028] = 8'b00000000;
dat[2029] = 8'b00000000;
dat[2030] = 8'b00000000;
dat[2031] = 8'b00000000;
dat[2032] = 8'b00000000;
dat[2033] = 8'b00000000;
dat[2034] = 8'b00000000;
dat[2035] = 8'b00000000;
dat[2036] = 8'b00000000;
dat[2037] = 8'b00000000;
dat[2038] = 8'b00000000;
dat[2039] = 8'b00000000;
dat[2040] = 8'b00000000;
dat[2041] = 8'b00000000;
dat[2042] = 8'b00000000;
dat[2043] = 8'b00000000;
dat[2044] = 8'b00000000;
dat[2045] = 8'b00000000;
dat[2046] = 8'b00000000;
dat[2047] = 8'b00000000;
dat[2048] = 8'b00000000;
dat[2049] = 8'b00000000;
dat[2050] = 8'b00000000;
dat[2051] = 8'b00000000;
dat[2052] = 8'b00000000;
dat[2053] = 8'b00000000;
dat[2054] = 8'b00000000;
dat[2055] = 8'b00000000;
dat[2056] = 8'b00000000;
dat[2057] = 8'b00000000;
dat[2058] = 8'b00000000;
dat[2059] = 8'b00000000;
dat[2060] = 8'b00000000;
dat[2061] = 8'b00000000;
dat[2062] = 8'b00000000;
dat[2063] = 8'b00000000;
dat[2064] = 8'b00000000;
dat[2065] = 8'b00000000;
dat[2066] = 8'b00000000;
dat[2067] = 8'b00000000;
dat[2068] = 8'b00000000;
dat[2069] = 8'b00000000;
dat[2070] = 8'b00000000;
dat[2071] = 8'b00000000;
dat[2072] = 8'b00000000;
dat[2073] = 8'b00000000;
dat[2074] = 8'b00000000;
dat[2075] = 8'b00000000;
dat[2076] = 8'b00000000;
dat[2077] = 8'b00000000;
dat[2078] = 8'b00000000;
dat[2079] = 8'b00000000;
dat[2080] = 8'b00000000;
dat[2081] = 8'b00000000;
dat[2082] = 8'b00000000;
dat[2083] = 8'b00000000;
dat[2084] = 8'b00000000;
dat[2085] = 8'b00000000;
dat[2086] = 8'b00000000;
dat[2087] = 8'b00000000;
dat[2088] = 8'b00000000;
dat[2089] = 8'b00000000;
dat[2090] = 8'b00000000;
dat[2091] = 8'b00000000;
dat[2092] = 8'b00000000;
dat[2093] = 8'b00000000;
dat[2094] = 8'b00000000;
dat[2095] = 8'b00000000;
dat[2096] = 8'b00000000;
dat[2097] = 8'b00000000;
dat[2098] = 8'b00000000;
dat[2099] = 8'b00000000;
dat[2100] = 8'b00000000;
dat[2101] = 8'b00000000;
dat[2102] = 8'b00000000;
dat[2103] = 8'b00000000;
dat[2104] = 8'b00000000;
dat[2105] = 8'b00000000;
dat[2106] = 8'b00000000;
dat[2107] = 8'b00000000;
dat[2108] = 8'b00000000;
dat[2109] = 8'b00000000;
dat[2110] = 8'b00000000;
dat[2111] = 8'b00000000;
dat[2112] = 8'b00000000;
dat[2113] = 8'b00000000;
dat[2114] = 8'b00000000;
dat[2115] = 8'b00000000;
dat[2116] = 8'b00000000;
dat[2117] = 8'b00000000;
dat[2118] = 8'b00000000;
dat[2119] = 8'b00000000;
dat[2120] = 8'b00000000;
dat[2121] = 8'b00000000;
dat[2122] = 8'b00000000;
dat[2123] = 8'b00000000;
dat[2124] = 8'b00000000;
dat[2125] = 8'b00000000;
dat[2126] = 8'b00000000;
dat[2127] = 8'b00000000;
dat[2128] = 8'b00000000;
dat[2129] = 8'b00000000;
dat[2130] = 8'b00000000;
dat[2131] = 8'b00000000;
dat[2132] = 8'b00000000;
dat[2133] = 8'b00000000;
dat[2134] = 8'b00000000;
dat[2135] = 8'b00000000;
dat[2136] = 8'b00000000;
dat[2137] = 8'b00000000;
dat[2138] = 8'b00000000;
dat[2139] = 8'b00000000;
dat[2140] = 8'b00000000;
dat[2141] = 8'b00000000;
dat[2142] = 8'b00000000;
dat[2143] = 8'b00000000;
dat[2144] = 8'b00000000;
dat[2145] = 8'b00000000;
dat[2146] = 8'b00000000;
dat[2147] = 8'b00000000;
dat[2148] = 8'b00000000;
dat[2149] = 8'b00000000;
dat[2150] = 8'b00000000;
dat[2151] = 8'b00000000;
dat[2152] = 8'b00000000;
dat[2153] = 8'b00000000;
dat[2154] = 8'b00000000;
dat[2155] = 8'b00000000;
dat[2156] = 8'b00000000;
dat[2157] = 8'b00000000;
dat[2158] = 8'b00000000;
dat[2159] = 8'b00000000;
dat[2160] = 8'b00000000;
dat[2161] = 8'b00000000;
dat[2162] = 8'b00000000;
dat[2163] = 8'b00000000;
dat[2164] = 8'b00000000;
dat[2165] = 8'b00000000;
dat[2166] = 8'b00000000;
dat[2167] = 8'b00000000;
dat[2168] = 8'b00000000;
dat[2169] = 8'b00000000;
dat[2170] = 8'b00000000;
dat[2171] = 8'b00000000;
dat[2172] = 8'b00000000;
dat[2173] = 8'b00000000;
dat[2174] = 8'b00000000;
dat[2175] = 8'b00000000;
dat[2176] = 8'b00000000;
dat[2177] = 8'b00000000;
dat[2178] = 8'b00000000;
dat[2179] = 8'b00000000;
dat[2180] = 8'b00000000;
dat[2181] = 8'b00000000;
dat[2182] = 8'b00000000;
dat[2183] = 8'b00000000;
dat[2184] = 8'b00000000;
dat[2185] = 8'b00000000;
dat[2186] = 8'b00000000;
dat[2187] = 8'b00000000;
dat[2188] = 8'b00000000;
dat[2189] = 8'b00000000;
dat[2190] = 8'b00000000;
dat[2191] = 8'b00000000;
dat[2192] = 8'b00000000;
dat[2193] = 8'b00000000;
dat[2194] = 8'b00000000;
dat[2195] = 8'b00000000;
dat[2196] = 8'b00000000;
dat[2197] = 8'b00000000;
dat[2198] = 8'b00000000;
dat[2199] = 8'b00000000;
dat[2200] = 8'b00000000;
dat[2201] = 8'b00000000;
dat[2202] = 8'b00000000;
dat[2203] = 8'b00000000;
dat[2204] = 8'b00000000;
dat[2205] = 8'b00000000;
dat[2206] = 8'b00000000;
dat[2207] = 8'b00000000;
dat[2208] = 8'b00000000;
dat[2209] = 8'b00000000;
dat[2210] = 8'b00000000;
dat[2211] = 8'b00000000;
dat[2212] = 8'b00000000;
dat[2213] = 8'b00000000;
dat[2214] = 8'b00000000;
dat[2215] = 8'b00000000;
dat[2216] = 8'b00000000;
dat[2217] = 8'b00000000;
dat[2218] = 8'b00000000;
dat[2219] = 8'b00000000;
dat[2220] = 8'b00000000;
dat[2221] = 8'b00000000;
dat[2222] = 8'b00000000;
dat[2223] = 8'b00000000;
dat[2224] = 8'b00000000;
dat[2225] = 8'b00000000;
dat[2226] = 8'b00000000;
dat[2227] = 8'b00000000;
dat[2228] = 8'b00000000;
dat[2229] = 8'b00000000;
dat[2230] = 8'b00000000;
dat[2231] = 8'b00000000;
dat[2232] = 8'b00000000;
dat[2233] = 8'b00000000;
dat[2234] = 8'b00000000;
dat[2235] = 8'b00000000;
dat[2236] = 8'b00000000;
dat[2237] = 8'b00000000;
dat[2238] = 8'b00000000;
dat[2239] = 8'b00000000;
dat[2240] = 8'b00000000;
dat[2241] = 8'b00000000;
dat[2242] = 8'b00000000;
dat[2243] = 8'b00000000;
dat[2244] = 8'b00000000;
dat[2245] = 8'b00000000;
dat[2246] = 8'b00000000;
dat[2247] = 8'b00000000;
dat[2248] = 8'b00000000;
dat[2249] = 8'b00000000;
dat[2250] = 8'b00000000;
dat[2251] = 8'b00000000;
dat[2252] = 8'b00000000;
dat[2253] = 8'b00000000;
dat[2254] = 8'b00000000;
dat[2255] = 8'b00000000;
dat[2256] = 8'b00000000;
dat[2257] = 8'b00000000;
dat[2258] = 8'b00000000;
dat[2259] = 8'b00000000;
dat[2260] = 8'b00000000;
dat[2261] = 8'b00000000;
dat[2262] = 8'b00000000;
dat[2263] = 8'b00000000;
dat[2264] = 8'b00000000;
dat[2265] = 8'b00000000;
dat[2266] = 8'b00000000;
dat[2267] = 8'b00000000;
dat[2268] = 8'b00000000;
dat[2269] = 8'b00000000;
dat[2270] = 8'b00000000;
dat[2271] = 8'b00000000;
dat[2272] = 8'b00000000;
dat[2273] = 8'b00000000;
dat[2274] = 8'b00000000;
dat[2275] = 8'b00000000;
dat[2276] = 8'b00000000;
dat[2277] = 8'b00000000;
dat[2278] = 8'b00000000;
dat[2279] = 8'b00000000;
dat[2280] = 8'b00000000;
dat[2281] = 8'b00000000;
dat[2282] = 8'b00000000;
dat[2283] = 8'b00000000;
dat[2284] = 8'b00000000;
dat[2285] = 8'b00000000;
dat[2286] = 8'b00000000;
dat[2287] = 8'b00000000;
dat[2288] = 8'b00000000;
dat[2289] = 8'b00000000;
dat[2290] = 8'b00000000;
dat[2291] = 8'b00000000;
dat[2292] = 8'b00000000;
dat[2293] = 8'b00000000;
dat[2294] = 8'b00000000;
dat[2295] = 8'b00000000;
dat[2296] = 8'b00000000;
dat[2297] = 8'b00000000;
dat[2298] = 8'b00000000;
dat[2299] = 8'b00000000;
dat[2300] = 8'b00000000;
dat[2301] = 8'b00000000;
dat[2302] = 8'b00000000;
dat[2303] = 8'b00000000;
dat[2304] = 8'b00000000;
dat[2305] = 8'b00000000;
dat[2306] = 8'b00000000;
dat[2307] = 8'b00000000;
dat[2308] = 8'b00000000;
dat[2309] = 8'b00000000;
dat[2310] = 8'b00000000;
dat[2311] = 8'b00000000;
dat[2312] = 8'b00000000;
dat[2313] = 8'b00000000;
dat[2314] = 8'b00000000;
dat[2315] = 8'b00000000;
dat[2316] = 8'b00000000;
dat[2317] = 8'b00000000;
dat[2318] = 8'b00000000;
dat[2319] = 8'b00000000;
dat[2320] = 8'b00000000;
dat[2321] = 8'b00000000;
dat[2322] = 8'b00000000;
dat[2323] = 8'b00000000;
dat[2324] = 8'b00000000;
dat[2325] = 8'b00000000;
dat[2326] = 8'b00000000;
dat[2327] = 8'b00000000;
dat[2328] = 8'b00000000;
dat[2329] = 8'b00000000;
dat[2330] = 8'b00000000;
dat[2331] = 8'b00000000;
dat[2332] = 8'b00000000;
dat[2333] = 8'b00000000;
dat[2334] = 8'b00000000;
dat[2335] = 8'b00000000;
dat[2336] = 8'b00000000;
dat[2337] = 8'b00000000;
dat[2338] = 8'b00000000;
dat[2339] = 8'b00000000;
dat[2340] = 8'b00000000;
dat[2341] = 8'b00000000;
dat[2342] = 8'b00000000;
dat[2343] = 8'b00000000;
dat[2344] = 8'b00000000;
dat[2345] = 8'b00000000;
dat[2346] = 8'b00000000;
dat[2347] = 8'b00000000;
dat[2348] = 8'b00000000;
dat[2349] = 8'b00000000;
dat[2350] = 8'b00000000;
dat[2351] = 8'b00000000;
dat[2352] = 8'b00000000;
dat[2353] = 8'b00000000;
dat[2354] = 8'b00000000;
dat[2355] = 8'b00000000;
dat[2356] = 8'b00000000;
dat[2357] = 8'b00000000;
dat[2358] = 8'b00000000;
dat[2359] = 8'b00000000;
dat[2360] = 8'b00000000;
dat[2361] = 8'b00000000;
dat[2362] = 8'b00000000;
dat[2363] = 8'b00000000;
dat[2364] = 8'b00000000;
dat[2365] = 8'b00000000;
dat[2366] = 8'b00000000;
dat[2367] = 8'b00000000;
dat[2368] = 8'b00000000;
dat[2369] = 8'b00000000;
dat[2370] = 8'b00000000;
dat[2371] = 8'b00000000;
dat[2372] = 8'b00000000;
dat[2373] = 8'b00000000;
dat[2374] = 8'b00000000;
dat[2375] = 8'b00000000;
dat[2376] = 8'b00000000;
dat[2377] = 8'b00000000;
dat[2378] = 8'b00000000;
dat[2379] = 8'b00000000;
dat[2380] = 8'b00000000;
dat[2381] = 8'b00000000;
dat[2382] = 8'b00000000;
dat[2383] = 8'b00000000;
dat[2384] = 8'b00000000;
dat[2385] = 8'b00000000;
dat[2386] = 8'b00000000;
dat[2387] = 8'b00000000;
dat[2388] = 8'b00000000;
dat[2389] = 8'b00000000;
dat[2390] = 8'b00000000;
dat[2391] = 8'b00000000;
dat[2392] = 8'b00000000;
dat[2393] = 8'b00000000;
dat[2394] = 8'b00000000;
dat[2395] = 8'b00000000;
dat[2396] = 8'b00000000;
dat[2397] = 8'b00000000;
dat[2398] = 8'b00000000;
dat[2399] = 8'b00000000;
dat[2400] = 8'b00000000;
dat[2401] = 8'b00000000;
dat[2402] = 8'b00000000;
dat[2403] = 8'b00000000;
dat[2404] = 8'b00000000;
dat[2405] = 8'b00000000;
dat[2406] = 8'b00000000;
dat[2407] = 8'b00000000;
dat[2408] = 8'b00000000;
dat[2409] = 8'b00000000;
dat[2410] = 8'b00000000;
dat[2411] = 8'b00000000;
dat[2412] = 8'b00000000;
dat[2413] = 8'b00000000;
dat[2414] = 8'b00000000;
dat[2415] = 8'b00000000;
dat[2416] = 8'b00000000;
dat[2417] = 8'b00000000;
dat[2418] = 8'b00000000;
dat[2419] = 8'b00000000;
dat[2420] = 8'b00000000;
dat[2421] = 8'b00000000;
dat[2422] = 8'b00000000;
dat[2423] = 8'b00000000;
dat[2424] = 8'b00000000;
dat[2425] = 8'b00000000;
dat[2426] = 8'b00000000;
dat[2427] = 8'b00000000;
dat[2428] = 8'b00000000;
dat[2429] = 8'b00000000;
dat[2430] = 8'b00000000;
dat[2431] = 8'b00000000;
dat[2432] = 8'b00000000;
dat[2433] = 8'b00000000;
dat[2434] = 8'b00000000;
dat[2435] = 8'b00000000;
dat[2436] = 8'b00000000;
dat[2437] = 8'b00000000;
dat[2438] = 8'b00000000;
dat[2439] = 8'b00000000;
dat[2440] = 8'b00000000;
dat[2441] = 8'b00000000;
dat[2442] = 8'b00000000;
dat[2443] = 8'b00000000;
dat[2444] = 8'b00000000;
dat[2445] = 8'b00000000;
dat[2446] = 8'b00000000;
dat[2447] = 8'b00000000;
dat[2448] = 8'b00000000;
dat[2449] = 8'b00000000;
dat[2450] = 8'b00000000;
dat[2451] = 8'b00000000;
dat[2452] = 8'b00000000;
dat[2453] = 8'b00000000;
dat[2454] = 8'b00000000;
dat[2455] = 8'b00000000;
dat[2456] = 8'b00000000;
dat[2457] = 8'b00000000;
dat[2458] = 8'b00000000;
dat[2459] = 8'b00000000;
dat[2460] = 8'b00000000;
dat[2461] = 8'b00000000;
dat[2462] = 8'b00000000;
dat[2463] = 8'b00000000;
dat[2464] = 8'b00000000;
dat[2465] = 8'b00000000;
dat[2466] = 8'b00000000;
dat[2467] = 8'b00000000;
dat[2468] = 8'b00000000;
dat[2469] = 8'b00000000;
dat[2470] = 8'b00000000;
dat[2471] = 8'b00000000;
dat[2472] = 8'b00000000;
dat[2473] = 8'b00000000;
dat[2474] = 8'b00000000;
dat[2475] = 8'b00000000;
dat[2476] = 8'b00000000;
dat[2477] = 8'b00000000;
dat[2478] = 8'b00000000;
dat[2479] = 8'b00000000;
dat[2480] = 8'b00000000;
dat[2481] = 8'b00000000;
dat[2482] = 8'b00000000;
dat[2483] = 8'b00000000;
dat[2484] = 8'b00000000;
dat[2485] = 8'b00000000;
dat[2486] = 8'b00000000;
dat[2487] = 8'b00000000;
dat[2488] = 8'b00000000;
dat[2489] = 8'b00000000;
dat[2490] = 8'b00000000;
dat[2491] = 8'b00000000;
dat[2492] = 8'b00000000;
dat[2493] = 8'b00000000;
dat[2494] = 8'b00000000;
dat[2495] = 8'b00000000;
dat[2496] = 8'b00000000;
dat[2497] = 8'b00000000;
dat[2498] = 8'b00000000;
dat[2499] = 8'b00000000;
dat[2500] = 8'b00000000;
dat[2501] = 8'b00000000;
dat[2502] = 8'b00000000;
dat[2503] = 8'b00000000;
dat[2504] = 8'b00000000;
dat[2505] = 8'b00000000;
dat[2506] = 8'b00000000;
dat[2507] = 8'b00000000;
dat[2508] = 8'b00000000;
dat[2509] = 8'b00000000;
dat[2510] = 8'b00000000;
dat[2511] = 8'b00000000;
dat[2512] = 8'b00000000;
dat[2513] = 8'b00000000;
dat[2514] = 8'b00000000;
dat[2515] = 8'b00000000;
dat[2516] = 8'b00000000;
dat[2517] = 8'b00000000;
dat[2518] = 8'b00000000;
dat[2519] = 8'b00000000;
dat[2520] = 8'b00000000;
dat[2521] = 8'b00000000;
dat[2522] = 8'b00000000;
dat[2523] = 8'b00000000;
dat[2524] = 8'b00000000;
dat[2525] = 8'b00000000;
dat[2526] = 8'b00000000;
dat[2527] = 8'b00000000;
dat[2528] = 8'b00000000;
dat[2529] = 8'b00000000;
dat[2530] = 8'b00000000;
dat[2531] = 8'b00000000;
dat[2532] = 8'b00000000;
dat[2533] = 8'b00000000;
dat[2534] = 8'b00000000;
dat[2535] = 8'b00000000;
dat[2536] = 8'b00000000;
dat[2537] = 8'b00000000;
dat[2538] = 8'b00000000;
dat[2539] = 8'b00000000;
dat[2540] = 8'b00000000;
dat[2541] = 8'b00000000;
dat[2542] = 8'b00000000;
dat[2543] = 8'b00000000;
dat[2544] = 8'b00000000;
dat[2545] = 8'b00000000;
dat[2546] = 8'b00000000;
dat[2547] = 8'b00000000;
dat[2548] = 8'b00000000;
dat[2549] = 8'b00000000;
dat[2550] = 8'b00000000;
dat[2551] = 8'b00000000;
dat[2552] = 8'b00000000;
dat[2553] = 8'b00000000;
dat[2554] = 8'b00000000;
dat[2555] = 8'b00000000;
dat[2556] = 8'b00000000;
dat[2557] = 8'b00000000;
dat[2558] = 8'b00000000;
dat[2559] = 8'b00000000;
dat[2560] = 8'b00000000;
dat[2561] = 8'b00000000;
dat[2562] = 8'b00000000;
dat[2563] = 8'b00000000;
dat[2564] = 8'b00000000;
dat[2565] = 8'b00000000;
dat[2566] = 8'b00000000;
dat[2567] = 8'b00000000;
dat[2568] = 8'b00000000;
dat[2569] = 8'b00000000;
dat[2570] = 8'b00000000;
dat[2571] = 8'b00000000;
dat[2572] = 8'b00000000;
dat[2573] = 8'b00000000;
dat[2574] = 8'b00000000;
dat[2575] = 8'b00000000;
dat[2576] = 8'b00000000;
dat[2577] = 8'b00000000;
dat[2578] = 8'b00000000;
dat[2579] = 8'b00000000;
dat[2580] = 8'b00000000;
dat[2581] = 8'b00000000;
dat[2582] = 8'b00000000;
dat[2583] = 8'b00000000;
dat[2584] = 8'b00000000;
dat[2585] = 8'b00000000;
dat[2586] = 8'b00000000;
dat[2587] = 8'b00000000;
dat[2588] = 8'b00000000;
dat[2589] = 8'b00000000;
dat[2590] = 8'b00000000;
dat[2591] = 8'b00000000;
dat[2592] = 8'b00000000;
dat[2593] = 8'b00000000;
dat[2594] = 8'b00000000;
dat[2595] = 8'b00000000;
dat[2596] = 8'b00000000;
dat[2597] = 8'b00000000;
dat[2598] = 8'b00000000;
dat[2599] = 8'b00000000;
dat[2600] = 8'b00000000;
dat[2601] = 8'b00000000;
dat[2602] = 8'b00000000;
dat[2603] = 8'b00000000;
dat[2604] = 8'b00000000;
dat[2605] = 8'b00000000;
dat[2606] = 8'b00000000;
dat[2607] = 8'b00000000;
dat[2608] = 8'b00000000;
dat[2609] = 8'b00000000;
dat[2610] = 8'b00000000;
dat[2611] = 8'b00000000;
dat[2612] = 8'b00000000;
dat[2613] = 8'b00000000;
dat[2614] = 8'b00000000;
dat[2615] = 8'b00000000;
dat[2616] = 8'b00000000;
dat[2617] = 8'b00000000;
dat[2618] = 8'b00000000;
dat[2619] = 8'b00000000;
dat[2620] = 8'b00000000;
dat[2621] = 8'b00000000;
dat[2622] = 8'b00000000;
dat[2623] = 8'b00000000;
dat[2624] = 8'b00000000;
dat[2625] = 8'b00000000;
dat[2626] = 8'b00000000;
dat[2627] = 8'b00000000;
dat[2628] = 8'b00000000;
dat[2629] = 8'b00000000;
dat[2630] = 8'b00000000;
dat[2631] = 8'b00000000;
dat[2632] = 8'b00000000;
dat[2633] = 8'b00000000;
dat[2634] = 8'b00000000;
dat[2635] = 8'b00000000;
dat[2636] = 8'b00000000;
dat[2637] = 8'b00000000;
dat[2638] = 8'b00000000;
dat[2639] = 8'b00000000;
dat[2640] = 8'b00000000;
dat[2641] = 8'b00000000;
dat[2642] = 8'b00000000;
dat[2643] = 8'b00000000;
dat[2644] = 8'b00000000;
dat[2645] = 8'b00000000;
dat[2646] = 8'b00000000;
dat[2647] = 8'b00000000;
dat[2648] = 8'b00000000;
dat[2649] = 8'b00000000;
dat[2650] = 8'b00000000;
dat[2651] = 8'b00000000;
dat[2652] = 8'b00000000;
dat[2653] = 8'b00000000;
dat[2654] = 8'b00000000;
dat[2655] = 8'b00000000;
dat[2656] = 8'b00000000;
dat[2657] = 8'b00000000;
dat[2658] = 8'b00000000;
dat[2659] = 8'b00000000;
dat[2660] = 8'b00000000;
dat[2661] = 8'b00000000;
dat[2662] = 8'b00000000;
dat[2663] = 8'b00000000;
dat[2664] = 8'b00000000;
dat[2665] = 8'b00000000;
dat[2666] = 8'b00000000;
dat[2667] = 8'b00000000;
dat[2668] = 8'b00000000;
dat[2669] = 8'b00000000;
dat[2670] = 8'b00000000;
dat[2671] = 8'b00000000;
dat[2672] = 8'b00000000;
dat[2673] = 8'b00000000;
dat[2674] = 8'b00000000;
dat[2675] = 8'b00000000;
dat[2676] = 8'b00000000;
dat[2677] = 8'b00000000;
dat[2678] = 8'b00000000;
dat[2679] = 8'b00000000;
dat[2680] = 8'b00000000;
dat[2681] = 8'b00000000;
dat[2682] = 8'b00000000;
dat[2683] = 8'b00000000;
dat[2684] = 8'b00000000;
dat[2685] = 8'b00000000;
dat[2686] = 8'b00000000;
dat[2687] = 8'b00000000;
dat[2688] = 8'b00000000;
dat[2689] = 8'b00000000;
dat[2690] = 8'b00000000;
dat[2691] = 8'b00000000;
dat[2692] = 8'b00000000;
dat[2693] = 8'b00000000;
dat[2694] = 8'b00000000;
dat[2695] = 8'b00000000;
dat[2696] = 8'b00000000;
dat[2697] = 8'b00000000;
dat[2698] = 8'b00000000;
dat[2699] = 8'b00000000;
dat[2700] = 8'b00000000;
dat[2701] = 8'b00000000;
dat[2702] = 8'b00000000;
dat[2703] = 8'b00000000;
dat[2704] = 8'b00000000;
dat[2705] = 8'b00000000;
dat[2706] = 8'b00000000;
dat[2707] = 8'b00000000;
dat[2708] = 8'b00000000;
dat[2709] = 8'b00000000;
dat[2710] = 8'b00000000;
dat[2711] = 8'b00000000;
dat[2712] = 8'b00000000;
dat[2713] = 8'b00000000;
dat[2714] = 8'b00000000;
dat[2715] = 8'b00000000;
dat[2716] = 8'b00000000;
dat[2717] = 8'b00000000;
dat[2718] = 8'b00000000;
dat[2719] = 8'b00000000;
dat[2720] = 8'b00000000;
dat[2721] = 8'b00000000;
dat[2722] = 8'b00000000;
dat[2723] = 8'b00000000;
dat[2724] = 8'b00000000;
dat[2725] = 8'b00000000;
dat[2726] = 8'b00000000;
dat[2727] = 8'b00000000;
dat[2728] = 8'b00000000;
dat[2729] = 8'b00000000;
dat[2730] = 8'b00000000;
dat[2731] = 8'b00000000;
dat[2732] = 8'b00000000;
dat[2733] = 8'b00000000;
dat[2734] = 8'b00000000;
dat[2735] = 8'b00000000;
dat[2736] = 8'b00000000;
dat[2737] = 8'b00000000;
dat[2738] = 8'b00000000;
dat[2739] = 8'b00000000;
dat[2740] = 8'b00000000;
dat[2741] = 8'b00000000;
dat[2742] = 8'b00000000;
dat[2743] = 8'b00000000;
dat[2744] = 8'b00000000;
dat[2745] = 8'b00000000;
dat[2746] = 8'b00000000;
dat[2747] = 8'b00000000;
dat[2748] = 8'b00000000;
dat[2749] = 8'b00000000;
dat[2750] = 8'b00000000;
dat[2751] = 8'b00000000;
dat[2752] = 8'b00000000;
dat[2753] = 8'b00000000;
dat[2754] = 8'b00000000;
dat[2755] = 8'b00000000;
dat[2756] = 8'b00000000;
dat[2757] = 8'b00000000;
dat[2758] = 8'b00000000;
dat[2759] = 8'b00000000;
dat[2760] = 8'b00000000;
dat[2761] = 8'b00000000;
dat[2762] = 8'b00000000;
dat[2763] = 8'b00000000;
dat[2764] = 8'b00000000;
dat[2765] = 8'b00000000;
dat[2766] = 8'b00000000;
dat[2767] = 8'b00000000;
dat[2768] = 8'b00000000;
dat[2769] = 8'b00000000;
dat[2770] = 8'b00000000;
dat[2771] = 8'b00000000;
dat[2772] = 8'b00000000;
dat[2773] = 8'b00000000;
dat[2774] = 8'b00000000;
dat[2775] = 8'b00000000;
dat[2776] = 8'b00000000;
dat[2777] = 8'b00000000;
dat[2778] = 8'b00000000;
dat[2779] = 8'b00000000;
dat[2780] = 8'b00000000;
dat[2781] = 8'b00000000;
dat[2782] = 8'b00000000;
dat[2783] = 8'b00000000;
dat[2784] = 8'b00000000;
dat[2785] = 8'b00000000;
dat[2786] = 8'b00000000;
dat[2787] = 8'b00000000;
dat[2788] = 8'b00000000;
dat[2789] = 8'b00000000;
dat[2790] = 8'b00000000;
dat[2791] = 8'b00000000;
dat[2792] = 8'b00000000;
dat[2793] = 8'b00000000;
dat[2794] = 8'b00000000;
dat[2795] = 8'b00000000;
dat[2796] = 8'b00000000;
dat[2797] = 8'b00000000;
dat[2798] = 8'b00000000;
dat[2799] = 8'b00000000;
dat[2800] = 8'b00000000;
dat[2801] = 8'b00000000;
dat[2802] = 8'b00000000;
dat[2803] = 8'b00000000;
dat[2804] = 8'b00000000;
dat[2805] = 8'b00000000;
dat[2806] = 8'b00000000;
dat[2807] = 8'b00000000;
dat[2808] = 8'b00000000;
dat[2809] = 8'b00000000;
dat[2810] = 8'b00000000;
dat[2811] = 8'b00000000;
dat[2812] = 8'b00000000;
dat[2813] = 8'b00000000;
dat[2814] = 8'b00000000;
dat[2815] = 8'b00000000;
dat[2816] = 8'b00000000;
dat[2817] = 8'b00000000;
dat[2818] = 8'b00000000;
dat[2819] = 8'b00000000;
dat[2820] = 8'b00000000;
dat[2821] = 8'b00000000;
dat[2822] = 8'b00000000;
dat[2823] = 8'b00000000;
dat[2824] = 8'b00000000;
dat[2825] = 8'b00000000;
dat[2826] = 8'b00000000;
dat[2827] = 8'b00000000;
dat[2828] = 8'b00000000;
dat[2829] = 8'b00000000;
dat[2830] = 8'b00000000;
dat[2831] = 8'b00000000;
dat[2832] = 8'b00000000;
dat[2833] = 8'b00000000;
dat[2834] = 8'b00000000;
dat[2835] = 8'b00000000;
dat[2836] = 8'b00000000;
dat[2837] = 8'b00000000;
dat[2838] = 8'b00000000;
dat[2839] = 8'b00000000;
dat[2840] = 8'b00000000;
dat[2841] = 8'b00000000;
dat[2842] = 8'b00000000;
dat[2843] = 8'b00000000;
dat[2844] = 8'b00000000;
dat[2845] = 8'b00000000;
dat[2846] = 8'b00000000;
dat[2847] = 8'b00000000;
dat[2848] = 8'b00000000;
dat[2849] = 8'b00000000;
dat[2850] = 8'b00000000;
dat[2851] = 8'b00000000;
dat[2852] = 8'b00000000;
dat[2853] = 8'b00000000;
dat[2854] = 8'b00000000;
dat[2855] = 8'b00000000;
dat[2856] = 8'b00000000;
dat[2857] = 8'b00000000;
dat[2858] = 8'b00000000;
dat[2859] = 8'b00000000;
dat[2860] = 8'b00000000;
dat[2861] = 8'b00000000;
dat[2862] = 8'b00000000;
dat[2863] = 8'b00000000;
dat[2864] = 8'b00000000;
dat[2865] = 8'b00000000;
dat[2866] = 8'b00000000;
dat[2867] = 8'b00000000;
dat[2868] = 8'b00000000;
dat[2869] = 8'b00000000;
dat[2870] = 8'b00000000;
dat[2871] = 8'b00000000;
dat[2872] = 8'b00000000;
dat[2873] = 8'b00000000;
dat[2874] = 8'b00000000;
dat[2875] = 8'b00000000;
dat[2876] = 8'b00000000;
dat[2877] = 8'b00000000;
dat[2878] = 8'b00000000;
dat[2879] = 8'b00000000;
dat[2880] = 8'b00000000;
dat[2881] = 8'b00000000;
dat[2882] = 8'b00000000;
dat[2883] = 8'b00000000;
dat[2884] = 8'b00000000;
dat[2885] = 8'b00000000;
dat[2886] = 8'b00000000;
dat[2887] = 8'b00000000;
dat[2888] = 8'b00000000;
dat[2889] = 8'b00000000;
dat[2890] = 8'b00000000;
dat[2891] = 8'b00000000;
dat[2892] = 8'b00000000;
dat[2893] = 8'b00000000;
dat[2894] = 8'b00000000;
dat[2895] = 8'b00000000;
dat[2896] = 8'b00000000;
dat[2897] = 8'b00000000;
dat[2898] = 8'b00000000;
dat[2899] = 8'b00000000;
dat[2900] = 8'b00000000;
dat[2901] = 8'b00000000;
dat[2902] = 8'b00000000;
dat[2903] = 8'b00000000;
dat[2904] = 8'b00000000;
dat[2905] = 8'b00000000;
dat[2906] = 8'b00000000;
dat[2907] = 8'b00000000;
dat[2908] = 8'b00000000;
dat[2909] = 8'b00000000;
dat[2910] = 8'b00000000;
dat[2911] = 8'b00000000;
dat[2912] = 8'b00000000;
dat[2913] = 8'b00000000;
dat[2914] = 8'b00000000;
dat[2915] = 8'b00000000;
dat[2916] = 8'b00000000;
dat[2917] = 8'b00000000;
dat[2918] = 8'b00000000;
dat[2919] = 8'b00000000;
dat[2920] = 8'b00000000;
dat[2921] = 8'b00000000;
dat[2922] = 8'b00000000;
dat[2923] = 8'b00000000;
dat[2924] = 8'b00000000;
dat[2925] = 8'b00000000;
dat[2926] = 8'b00000000;
dat[2927] = 8'b00000000;
dat[2928] = 8'b00000000;
dat[2929] = 8'b00000000;
dat[2930] = 8'b00000000;
dat[2931] = 8'b00000000;
dat[2932] = 8'b00000000;
dat[2933] = 8'b00000000;
dat[2934] = 8'b00000000;
dat[2935] = 8'b00000000;
dat[2936] = 8'b00000000;
dat[2937] = 8'b00000000;
dat[2938] = 8'b00000000;
dat[2939] = 8'b00000000;
dat[2940] = 8'b00000000;
dat[2941] = 8'b00000000;
dat[2942] = 8'b00000000;
dat[2943] = 8'b00000000;
dat[2944] = 8'b00000000;
dat[2945] = 8'b00000000;
dat[2946] = 8'b00000000;
dat[2947] = 8'b00000000;
dat[2948] = 8'b00000000;
dat[2949] = 8'b00000000;
dat[2950] = 8'b00000000;
dat[2951] = 8'b00000000;
dat[2952] = 8'b00000000;
dat[2953] = 8'b00000000;
dat[2954] = 8'b00000000;
dat[2955] = 8'b00000000;
dat[2956] = 8'b00000000;
dat[2957] = 8'b00000000;
dat[2958] = 8'b00000000;
dat[2959] = 8'b00000000;
dat[2960] = 8'b00000000;
dat[2961] = 8'b00000000;
dat[2962] = 8'b00000000;
dat[2963] = 8'b00000000;
dat[2964] = 8'b00000000;
dat[2965] = 8'b00000000;
dat[2966] = 8'b00000000;
dat[2967] = 8'b00000000;
dat[2968] = 8'b00000000;
dat[2969] = 8'b00000000;
dat[2970] = 8'b00000000;
dat[2971] = 8'b00000000;
dat[2972] = 8'b00000000;
dat[2973] = 8'b00000000;
dat[2974] = 8'b00000000;
dat[2975] = 8'b00000000;
dat[2976] = 8'b00000000;
dat[2977] = 8'b00000000;
dat[2978] = 8'b00000000;
dat[2979] = 8'b00000000;
dat[2980] = 8'b00000000;
dat[2981] = 8'b00000000;
dat[2982] = 8'b00000000;
dat[2983] = 8'b00000000;
dat[2984] = 8'b00000000;
dat[2985] = 8'b00000000;
dat[2986] = 8'b00000000;
dat[2987] = 8'b00000000;
dat[2988] = 8'b00000000;
dat[2989] = 8'b00000000;
dat[2990] = 8'b00000000;
dat[2991] = 8'b00000000;
dat[2992] = 8'b00000000;
dat[2993] = 8'b00000000;
dat[2994] = 8'b00000000;
dat[2995] = 8'b00000000;
dat[2996] = 8'b00000000;
dat[2997] = 8'b00000000;
dat[2998] = 8'b00000000;
dat[2999] = 8'b00000000;
dat[3000] = 8'b00000000;
dat[3001] = 8'b00000000;
dat[3002] = 8'b00000000;
dat[3003] = 8'b00000000;
dat[3004] = 8'b00000000;
dat[3005] = 8'b00000000;
dat[3006] = 8'b00000000;
dat[3007] = 8'b00000000;
dat[3008] = 8'b00000000;
dat[3009] = 8'b00000000;
dat[3010] = 8'b00000000;
dat[3011] = 8'b00000000;
dat[3012] = 8'b00000000;
dat[3013] = 8'b00000000;
dat[3014] = 8'b00000000;
dat[3015] = 8'b00000000;
dat[3016] = 8'b00000000;
dat[3017] = 8'b00000000;
dat[3018] = 8'b00000000;
dat[3019] = 8'b00000000;
dat[3020] = 8'b00000000;
dat[3021] = 8'b00000000;
dat[3022] = 8'b00000000;
dat[3023] = 8'b00000000;
dat[3024] = 8'b00000000;
dat[3025] = 8'b00000000;
dat[3026] = 8'b00000000;
dat[3027] = 8'b00000000;
dat[3028] = 8'b00000000;
dat[3029] = 8'b00000000;
dat[3030] = 8'b00000000;
dat[3031] = 8'b00000000;
dat[3032] = 8'b00000000;
dat[3033] = 8'b00000000;
dat[3034] = 8'b00000000;
dat[3035] = 8'b00000000;
dat[3036] = 8'b00000000;
dat[3037] = 8'b00000000;
dat[3038] = 8'b00000000;
dat[3039] = 8'b00000000;
dat[3040] = 8'b00000000;
dat[3041] = 8'b00000000;
dat[3042] = 8'b00000000;
dat[3043] = 8'b00000000;
dat[3044] = 8'b00000000;
dat[3045] = 8'b00000000;
dat[3046] = 8'b00000000;
dat[3047] = 8'b00000000;
dat[3048] = 8'b00000000;
dat[3049] = 8'b00000000;
dat[3050] = 8'b00000000;
dat[3051] = 8'b00000000;
dat[3052] = 8'b00000000;
dat[3053] = 8'b00000000;
dat[3054] = 8'b00000000;
dat[3055] = 8'b00000000;
dat[3056] = 8'b00000000;
dat[3057] = 8'b00000000;
dat[3058] = 8'b00000000;
dat[3059] = 8'b00000000;
dat[3060] = 8'b00000000;
dat[3061] = 8'b00000000;
dat[3062] = 8'b00000000;
dat[3063] = 8'b00000000;
dat[3064] = 8'b00000000;
dat[3065] = 8'b00000000;
dat[3066] = 8'b00000000;
dat[3067] = 8'b00000000;
dat[3068] = 8'b00000000;
dat[3069] = 8'b00000000;
dat[3070] = 8'b00000000;
dat[3071] = 8'b00000000;
dat[3072] = 8'b00000000;
dat[3073] = 8'b00000000;
dat[3074] = 8'b00000000;
dat[3075] = 8'b00000000;
dat[3076] = 8'b00000000;
dat[3077] = 8'b00000000;
dat[3078] = 8'b00000000;
dat[3079] = 8'b00000000;
dat[3080] = 8'b00000000;
dat[3081] = 8'b00000000;
dat[3082] = 8'b00000000;
dat[3083] = 8'b00000000;
dat[3084] = 8'b00000000;
dat[3085] = 8'b00000000;
dat[3086] = 8'b00000000;
dat[3087] = 8'b00000000;
dat[3088] = 8'b00000000;
dat[3089] = 8'b00000000;
dat[3090] = 8'b00000000;
dat[3091] = 8'b00000000;
dat[3092] = 8'b00000000;
dat[3093] = 8'b00000000;
dat[3094] = 8'b00000000;
dat[3095] = 8'b00000000;
dat[3096] = 8'b00000000;
dat[3097] = 8'b00000000;
dat[3098] = 8'b00000000;
dat[3099] = 8'b00000000;
dat[3100] = 8'b00000000;
dat[3101] = 8'b00000000;
dat[3102] = 8'b00000000;
dat[3103] = 8'b00000000;
dat[3104] = 8'b00000000;
dat[3105] = 8'b00000000;
dat[3106] = 8'b00000000;
dat[3107] = 8'b00000000;
dat[3108] = 8'b00000000;
dat[3109] = 8'b00000000;
dat[3110] = 8'b00000000;
dat[3111] = 8'b00000000;
dat[3112] = 8'b00000000;
dat[3113] = 8'b00000000;
dat[3114] = 8'b00000000;
dat[3115] = 8'b00000000;
dat[3116] = 8'b00000000;
dat[3117] = 8'b00000000;
dat[3118] = 8'b00000000;
dat[3119] = 8'b00000000;
dat[3120] = 8'b00000000;
dat[3121] = 8'b00000000;
dat[3122] = 8'b00000000;
dat[3123] = 8'b00000000;
dat[3124] = 8'b00000000;
dat[3125] = 8'b00000000;
dat[3126] = 8'b00000000;
dat[3127] = 8'b00000000;
dat[3128] = 8'b00000000;
dat[3129] = 8'b00000000;
dat[3130] = 8'b00000000;
dat[3131] = 8'b00000000;
dat[3132] = 8'b00000000;
dat[3133] = 8'b00000000;
dat[3134] = 8'b00000000;
dat[3135] = 8'b00000000;
dat[3136] = 8'b00000000;
dat[3137] = 8'b00000000;
dat[3138] = 8'b00000000;
dat[3139] = 8'b00000000;
dat[3140] = 8'b00000000;
dat[3141] = 8'b00000000;
dat[3142] = 8'b00000000;
dat[3143] = 8'b00000000;
dat[3144] = 8'b00000000;
dat[3145] = 8'b00000000;
dat[3146] = 8'b00000000;
dat[3147] = 8'b00000000;
dat[3148] = 8'b00000000;
dat[3149] = 8'b00000000;
dat[3150] = 8'b00000000;
dat[3151] = 8'b00000000;
dat[3152] = 8'b00000000;
dat[3153] = 8'b00000000;
dat[3154] = 8'b00000000;
dat[3155] = 8'b00000000;
dat[3156] = 8'b00000000;
dat[3157] = 8'b00000000;
dat[3158] = 8'b00000000;
dat[3159] = 8'b00000000;
dat[3160] = 8'b00000000;
dat[3161] = 8'b00000000;
dat[3162] = 8'b00000000;
dat[3163] = 8'b00000000;
dat[3164] = 8'b00000000;
dat[3165] = 8'b00000000;
dat[3166] = 8'b00000000;
dat[3167] = 8'b00000000;
dat[3168] = 8'b00000000;
dat[3169] = 8'b00000000;
dat[3170] = 8'b00000000;
dat[3171] = 8'b00000000;
dat[3172] = 8'b00000000;
dat[3173] = 8'b00000000;
dat[3174] = 8'b00000000;
dat[3175] = 8'b00000000;
dat[3176] = 8'b00000000;
dat[3177] = 8'b00000000;
dat[3178] = 8'b00000000;
dat[3179] = 8'b00000000;
dat[3180] = 8'b00000000;
dat[3181] = 8'b00000000;
dat[3182] = 8'b00000000;
dat[3183] = 8'b00000000;
dat[3184] = 8'b00000000;
dat[3185] = 8'b00000000;
dat[3186] = 8'b00000000;
dat[3187] = 8'b00000000;
dat[3188] = 8'b00000000;
dat[3189] = 8'b00000000;
dat[3190] = 8'b00000000;
dat[3191] = 8'b00000000;
dat[3192] = 8'b00000000;
dat[3193] = 8'b00000000;
dat[3194] = 8'b00000000;
dat[3195] = 8'b00000000;
dat[3196] = 8'b00000000;
dat[3197] = 8'b00000000;
dat[3198] = 8'b00000000;
dat[3199] = 8'b00000000;
dat[3200] = 8'b00000000;
dat[3201] = 8'b00000000;
dat[3202] = 8'b00000000;
dat[3203] = 8'b00000000;
dat[3204] = 8'b00000000;
dat[3205] = 8'b00000000;
dat[3206] = 8'b00000000;
dat[3207] = 8'b00000000;
dat[3208] = 8'b00000000;
dat[3209] = 8'b00000000;
dat[3210] = 8'b00000000;
dat[3211] = 8'b00000000;
dat[3212] = 8'b00000000;
dat[3213] = 8'b00000000;
dat[3214] = 8'b00000000;
dat[3215] = 8'b00000000;
dat[3216] = 8'b00000000;
dat[3217] = 8'b00000000;
dat[3218] = 8'b00000000;
dat[3219] = 8'b00000000;
dat[3220] = 8'b00000000;
dat[3221] = 8'b00000000;
dat[3222] = 8'b00000000;
dat[3223] = 8'b00000000;
dat[3224] = 8'b00000000;
dat[3225] = 8'b00000000;
dat[3226] = 8'b00000000;
dat[3227] = 8'b00000000;
dat[3228] = 8'b00000000;
dat[3229] = 8'b00000000;
dat[3230] = 8'b00000000;
dat[3231] = 8'b00000000;
dat[3232] = 8'b00000000;
dat[3233] = 8'b00000000;
dat[3234] = 8'b00000000;
dat[3235] = 8'b00000000;
dat[3236] = 8'b00000000;
dat[3237] = 8'b00000000;
dat[3238] = 8'b00000000;
dat[3239] = 8'b00000000;
dat[3240] = 8'b00000000;
dat[3241] = 8'b00000000;
dat[3242] = 8'b00000000;
dat[3243] = 8'b00000000;
dat[3244] = 8'b00000000;
dat[3245] = 8'b00000000;
dat[3246] = 8'b00000000;
dat[3247] = 8'b00000000;
dat[3248] = 8'b00000000;
dat[3249] = 8'b00000000;
dat[3250] = 8'b00000000;
dat[3251] = 8'b00000000;
dat[3252] = 8'b00000000;
dat[3253] = 8'b00000000;
dat[3254] = 8'b00000000;
dat[3255] = 8'b00000000;
dat[3256] = 8'b00000000;
dat[3257] = 8'b00000000;
dat[3258] = 8'b00000000;
dat[3259] = 8'b00000000;
dat[3260] = 8'b00000000;
dat[3261] = 8'b00000000;
dat[3262] = 8'b00000000;
dat[3263] = 8'b00000000;
dat[3264] = 8'b00000000;
dat[3265] = 8'b00000000;
dat[3266] = 8'b00000000;
dat[3267] = 8'b00000000;
dat[3268] = 8'b00000000;
dat[3269] = 8'b00000000;
dat[3270] = 8'b00000000;
dat[3271] = 8'b00000000;
dat[3272] = 8'b00000000;
dat[3273] = 8'b00000000;
dat[3274] = 8'b00000000;
dat[3275] = 8'b00000000;
dat[3276] = 8'b00000000;
dat[3277] = 8'b00000000;
dat[3278] = 8'b00000000;
dat[3279] = 8'b00000000;
dat[3280] = 8'b00000000;
dat[3281] = 8'b00000000;
dat[3282] = 8'b00000000;
dat[3283] = 8'b00000000;
dat[3284] = 8'b00000000;
dat[3285] = 8'b00000000;
dat[3286] = 8'b00000000;
dat[3287] = 8'b00000000;
dat[3288] = 8'b00000000;
dat[3289] = 8'b00000000;
dat[3290] = 8'b00000000;
dat[3291] = 8'b00000000;
dat[3292] = 8'b00000000;
dat[3293] = 8'b00000000;
dat[3294] = 8'b00000000;
dat[3295] = 8'b00000000;
dat[3296] = 8'b00000000;
dat[3297] = 8'b00000000;
dat[3298] = 8'b00000000;
dat[3299] = 8'b00000000;
dat[3300] = 8'b00000000;
dat[3301] = 8'b00000000;
dat[3302] = 8'b00000000;
dat[3303] = 8'b00000000;
dat[3304] = 8'b00000000;
dat[3305] = 8'b00000000;
dat[3306] = 8'b00000000;
dat[3307] = 8'b00000000;
dat[3308] = 8'b00000000;
dat[3309] = 8'b00000000;
dat[3310] = 8'b00000000;
dat[3311] = 8'b00000000;
dat[3312] = 8'b00000000;
dat[3313] = 8'b00000000;
dat[3314] = 8'b00000000;
dat[3315] = 8'b00000000;
dat[3316] = 8'b00000000;
dat[3317] = 8'b00000000;
dat[3318] = 8'b00000000;
dat[3319] = 8'b00000000;
dat[3320] = 8'b00000000;
dat[3321] = 8'b00000000;
dat[3322] = 8'b00000000;
dat[3323] = 8'b00000000;
dat[3324] = 8'b00000000;
dat[3325] = 8'b00000000;
dat[3326] = 8'b00000000;
dat[3327] = 8'b00000000;
dat[3328] = 8'b00000000;
dat[3329] = 8'b00000000;
dat[3330] = 8'b00000000;
dat[3331] = 8'b00000000;
dat[3332] = 8'b00000000;
dat[3333] = 8'b00000000;
dat[3334] = 8'b00000000;
dat[3335] = 8'b00000000;
dat[3336] = 8'b00000000;
dat[3337] = 8'b00000000;
dat[3338] = 8'b00000000;
dat[3339] = 8'b00000000;
dat[3340] = 8'b00000000;
dat[3341] = 8'b00000000;
dat[3342] = 8'b00000000;
dat[3343] = 8'b00000000;
dat[3344] = 8'b00000000;
dat[3345] = 8'b00000000;
dat[3346] = 8'b00000000;
dat[3347] = 8'b00000000;
dat[3348] = 8'b00000000;
dat[3349] = 8'b00000000;
dat[3350] = 8'b00000000;
dat[3351] = 8'b00000000;
dat[3352] = 8'b00000000;
dat[3353] = 8'b00000000;
dat[3354] = 8'b00000000;
dat[3355] = 8'b00000000;
dat[3356] = 8'b00000000;
dat[3357] = 8'b00000000;
dat[3358] = 8'b00000000;
dat[3359] = 8'b00000000;
dat[3360] = 8'b00000000;
dat[3361] = 8'b00000000;
dat[3362] = 8'b00000000;
dat[3363] = 8'b00000000;
dat[3364] = 8'b00000000;
dat[3365] = 8'b00000000;
dat[3366] = 8'b00000000;
dat[3367] = 8'b00000000;
dat[3368] = 8'b00000000;
dat[3369] = 8'b00000000;
dat[3370] = 8'b00000000;
dat[3371] = 8'b00000000;
dat[3372] = 8'b00000000;
dat[3373] = 8'b00000000;
dat[3374] = 8'b00000000;
dat[3375] = 8'b00000000;
dat[3376] = 8'b00000000;
dat[3377] = 8'b00000000;
dat[3378] = 8'b00000000;
dat[3379] = 8'b00000000;
dat[3380] = 8'b00000000;
dat[3381] = 8'b00000000;
dat[3382] = 8'b00000000;
dat[3383] = 8'b00000000;
dat[3384] = 8'b00000000;
dat[3385] = 8'b00000000;
dat[3386] = 8'b00000000;
dat[3387] = 8'b00000000;
dat[3388] = 8'b00000000;
dat[3389] = 8'b00000000;
dat[3390] = 8'b00000000;
dat[3391] = 8'b00000000;
dat[3392] = 8'b00000000;
dat[3393] = 8'b00000000;
dat[3394] = 8'b00000000;
dat[3395] = 8'b00000000;
dat[3396] = 8'b00000000;
dat[3397] = 8'b00000000;
dat[3398] = 8'b00000000;
dat[3399] = 8'b00000000;
dat[3400] = 8'b00000000;
dat[3401] = 8'b00000000;
dat[3402] = 8'b00000000;
dat[3403] = 8'b00000000;
dat[3404] = 8'b00000000;
dat[3405] = 8'b00000000;
dat[3406] = 8'b00000000;
dat[3407] = 8'b00000000;
dat[3408] = 8'b00000000;
dat[3409] = 8'b00000000;
dat[3410] = 8'b00000000;
dat[3411] = 8'b00000000;
dat[3412] = 8'b00000000;
dat[3413] = 8'b00000000;
dat[3414] = 8'b00000000;
dat[3415] = 8'b00000000;
dat[3416] = 8'b00000000;
dat[3417] = 8'b00000000;
dat[3418] = 8'b00000000;
dat[3419] = 8'b00000000;
dat[3420] = 8'b00000000;
dat[3421] = 8'b00000000;
dat[3422] = 8'b00000000;
dat[3423] = 8'b00000000;
dat[3424] = 8'b00000000;
dat[3425] = 8'b00000000;
dat[3426] = 8'b00000000;
dat[3427] = 8'b00000000;
dat[3428] = 8'b00000000;
dat[3429] = 8'b00000000;
dat[3430] = 8'b00000000;
dat[3431] = 8'b00000000;
dat[3432] = 8'b00000000;
dat[3433] = 8'b00000000;
dat[3434] = 8'b00000000;
dat[3435] = 8'b00000000;
dat[3436] = 8'b00000000;
dat[3437] = 8'b00000000;
dat[3438] = 8'b00000000;
dat[3439] = 8'b00000000;
dat[3440] = 8'b00000000;
dat[3441] = 8'b00000000;
dat[3442] = 8'b00000000;
dat[3443] = 8'b00000000;
dat[3444] = 8'b00000000;
dat[3445] = 8'b00000000;
dat[3446] = 8'b00000000;
dat[3447] = 8'b00000000;
dat[3448] = 8'b00000000;
dat[3449] = 8'b00000000;
dat[3450] = 8'b00000000;
dat[3451] = 8'b00000000;
dat[3452] = 8'b00000000;
dat[3453] = 8'b00000000;
dat[3454] = 8'b00000000;
dat[3455] = 8'b00000000;
dat[3456] = 8'b00000000;
dat[3457] = 8'b00000000;
dat[3458] = 8'b00000000;
dat[3459] = 8'b00000000;
dat[3460] = 8'b00000000;
dat[3461] = 8'b00000000;
dat[3462] = 8'b00000000;
dat[3463] = 8'b00000000;
dat[3464] = 8'b00000000;
dat[3465] = 8'b00000000;
dat[3466] = 8'b00000000;
dat[3467] = 8'b00000000;
dat[3468] = 8'b00000000;
dat[3469] = 8'b00000000;
dat[3470] = 8'b00000000;
dat[3471] = 8'b00000000;
dat[3472] = 8'b00000000;
dat[3473] = 8'b00000000;
dat[3474] = 8'b00000000;
dat[3475] = 8'b00000000;
dat[3476] = 8'b00000000;
dat[3477] = 8'b00000000;
dat[3478] = 8'b00000000;
dat[3479] = 8'b00000000;
dat[3480] = 8'b00000000;
dat[3481] = 8'b00000000;
dat[3482] = 8'b00000000;
dat[3483] = 8'b00000000;
dat[3484] = 8'b00000000;
dat[3485] = 8'b00000000;
dat[3486] = 8'b00000000;
dat[3487] = 8'b00000000;
dat[3488] = 8'b00000000;
dat[3489] = 8'b00000000;
dat[3490] = 8'b00000000;
dat[3491] = 8'b00000000;
dat[3492] = 8'b00000000;
dat[3493] = 8'b00000000;
dat[3494] = 8'b00000000;
dat[3495] = 8'b00000000;
dat[3496] = 8'b00000000;
dat[3497] = 8'b00000000;
dat[3498] = 8'b00000000;
dat[3499] = 8'b00000000;
dat[3500] = 8'b00000000;
dat[3501] = 8'b00000000;
dat[3502] = 8'b00000000;
dat[3503] = 8'b00000000;
dat[3504] = 8'b00000000;
dat[3505] = 8'b00000000;
dat[3506] = 8'b00000000;
dat[3507] = 8'b00000000;
dat[3508] = 8'b00000000;
dat[3509] = 8'b00000000;
dat[3510] = 8'b00000000;
dat[3511] = 8'b00000000;
dat[3512] = 8'b00000000;
dat[3513] = 8'b00000000;
dat[3514] = 8'b00000000;
dat[3515] = 8'b00000000;
dat[3516] = 8'b00000000;
dat[3517] = 8'b00000000;
dat[3518] = 8'b00000000;
dat[3519] = 8'b00000000;
dat[3520] = 8'b00000000;
dat[3521] = 8'b00000000;
dat[3522] = 8'b00000000;
dat[3523] = 8'b00000000;
dat[3524] = 8'b00000000;
dat[3525] = 8'b00000000;
dat[3526] = 8'b00000000;
dat[3527] = 8'b00000000;
dat[3528] = 8'b00000000;
dat[3529] = 8'b00000000;
dat[3530] = 8'b00000000;
dat[3531] = 8'b00000000;
dat[3532] = 8'b00000000;
dat[3533] = 8'b00000000;
dat[3534] = 8'b00000000;
dat[3535] = 8'b00000000;
dat[3536] = 8'b00000000;
dat[3537] = 8'b00000000;
dat[3538] = 8'b00000000;
dat[3539] = 8'b00000000;
dat[3540] = 8'b00000000;
dat[3541] = 8'b00000000;
dat[3542] = 8'b00000000;
dat[3543] = 8'b00000000;
dat[3544] = 8'b00000000;
dat[3545] = 8'b00000000;
dat[3546] = 8'b00000000;
dat[3547] = 8'b00000000;
dat[3548] = 8'b00000000;
dat[3549] = 8'b00000000;
dat[3550] = 8'b00000000;
dat[3551] = 8'b00000000;
dat[3552] = 8'b00000000;
dat[3553] = 8'b00000000;
dat[3554] = 8'b00000000;
dat[3555] = 8'b00000000;
dat[3556] = 8'b00000000;
dat[3557] = 8'b00000000;
dat[3558] = 8'b00000000;
dat[3559] = 8'b00000000;
dat[3560] = 8'b00000000;
dat[3561] = 8'b00000000;
dat[3562] = 8'b00000000;
dat[3563] = 8'b00000000;
dat[3564] = 8'b00000000;
dat[3565] = 8'b00000000;
dat[3566] = 8'b00000000;
dat[3567] = 8'b00000000;
dat[3568] = 8'b00000000;
dat[3569] = 8'b00000000;
dat[3570] = 8'b00000000;
dat[3571] = 8'b00000000;
dat[3572] = 8'b00000000;
dat[3573] = 8'b00000000;
dat[3574] = 8'b00000000;
dat[3575] = 8'b00000000;
dat[3576] = 8'b00000000;
dat[3577] = 8'b00000000;
dat[3578] = 8'b00000000;
dat[3579] = 8'b00000000;
dat[3580] = 8'b00000000;
dat[3581] = 8'b00000000;
dat[3582] = 8'b00000000;
dat[3583] = 8'b00000000;
dat[3584] = 8'b00000000;
dat[3585] = 8'b00000000;
dat[3586] = 8'b00000000;
dat[3587] = 8'b00000000;
dat[3588] = 8'b00000000;
dat[3589] = 8'b00000000;
dat[3590] = 8'b00000000;
dat[3591] = 8'b00000000;
dat[3592] = 8'b00000000;
dat[3593] = 8'b00000000;
dat[3594] = 8'b00000000;
dat[3595] = 8'b00000000;
dat[3596] = 8'b00000000;
dat[3597] = 8'b00000000;
dat[3598] = 8'b00000000;
dat[3599] = 8'b00000000;
dat[3600] = 8'b00000000;
dat[3601] = 8'b00000000;
dat[3602] = 8'b00000000;
dat[3603] = 8'b00000000;
dat[3604] = 8'b00000000;
dat[3605] = 8'b00000000;
dat[3606] = 8'b00000000;
dat[3607] = 8'b00000000;
dat[3608] = 8'b00000000;
dat[3609] = 8'b00000000;
dat[3610] = 8'b00000000;
dat[3611] = 8'b00000000;
dat[3612] = 8'b00000000;
dat[3613] = 8'b00000000;
dat[3614] = 8'b00000000;
dat[3615] = 8'b00000000;
dat[3616] = 8'b00000000;
dat[3617] = 8'b00000000;
dat[3618] = 8'b00000000;
dat[3619] = 8'b00000000;
dat[3620] = 8'b00000000;
dat[3621] = 8'b00000000;
dat[3622] = 8'b00000000;
dat[3623] = 8'b00000000;
dat[3624] = 8'b00000000;
dat[3625] = 8'b00000000;
dat[3626] = 8'b00000000;
dat[3627] = 8'b00000000;
dat[3628] = 8'b00000000;
dat[3629] = 8'b00000000;
dat[3630] = 8'b00000000;
dat[3631] = 8'b00000000;
dat[3632] = 8'b00000000;
dat[3633] = 8'b00000000;
dat[3634] = 8'b00000000;
dat[3635] = 8'b00000000;
dat[3636] = 8'b00000000;
dat[3637] = 8'b00000000;
dat[3638] = 8'b00000000;
dat[3639] = 8'b00000000;
dat[3640] = 8'b00000000;
dat[3641] = 8'b00000000;
dat[3642] = 8'b00000000;
dat[3643] = 8'b00000000;
dat[3644] = 8'b00000000;
dat[3645] = 8'b00000000;
dat[3646] = 8'b00000000;
dat[3647] = 8'b00000000;
dat[3648] = 8'b00000000;
dat[3649] = 8'b00000000;
dat[3650] = 8'b00000000;
dat[3651] = 8'b00000000;
dat[3652] = 8'b00000000;
dat[3653] = 8'b00000000;
dat[3654] = 8'b00000000;
dat[3655] = 8'b00000000;
dat[3656] = 8'b00000000;
dat[3657] = 8'b00000000;
dat[3658] = 8'b00000000;
dat[3659] = 8'b00000000;
dat[3660] = 8'b00000000;
dat[3661] = 8'b00000000;
dat[3662] = 8'b00000000;
dat[3663] = 8'b00000000;
dat[3664] = 8'b00000000;
dat[3665] = 8'b00000000;
dat[3666] = 8'b00000000;
dat[3667] = 8'b00000000;
dat[3668] = 8'b00000000;
dat[3669] = 8'b00000000;
dat[3670] = 8'b00000000;
dat[3671] = 8'b00000000;
dat[3672] = 8'b00000000;
dat[3673] = 8'b00000000;
dat[3674] = 8'b00000000;
dat[3675] = 8'b00000000;
dat[3676] = 8'b00000000;
dat[3677] = 8'b00000000;
dat[3678] = 8'b00000000;
dat[3679] = 8'b00000000;
dat[3680] = 8'b00000000;
dat[3681] = 8'b00000000;
dat[3682] = 8'b00000000;
dat[3683] = 8'b00000000;
dat[3684] = 8'b00000000;
dat[3685] = 8'b00000000;
dat[3686] = 8'b00000000;
dat[3687] = 8'b00000000;
dat[3688] = 8'b00000000;
dat[3689] = 8'b00000000;
dat[3690] = 8'b00000000;
dat[3691] = 8'b00000000;
dat[3692] = 8'b00000000;
dat[3693] = 8'b00000000;
dat[3694] = 8'b00000000;
dat[3695] = 8'b00000000;
dat[3696] = 8'b00000000;
dat[3697] = 8'b00000000;
dat[3698] = 8'b00000000;
dat[3699] = 8'b00000000;
dat[3700] = 8'b00000000;
dat[3701] = 8'b00000000;
dat[3702] = 8'b00000000;
dat[3703] = 8'b00000000;
dat[3704] = 8'b00000000;
dat[3705] = 8'b00000000;
dat[3706] = 8'b00000000;
dat[3707] = 8'b00000000;
dat[3708] = 8'b00000000;
dat[3709] = 8'b00000000;
dat[3710] = 8'b00000000;
dat[3711] = 8'b00000000;
dat[3712] = 8'b00000000;
dat[3713] = 8'b00000000;
dat[3714] = 8'b00000000;
dat[3715] = 8'b00000000;
dat[3716] = 8'b00000000;
dat[3717] = 8'b00000000;
dat[3718] = 8'b00000000;
dat[3719] = 8'b00000000;
dat[3720] = 8'b00000000;
dat[3721] = 8'b00000000;
dat[3722] = 8'b00000000;
dat[3723] = 8'b00000000;
dat[3724] = 8'b00000000;
dat[3725] = 8'b00000000;
dat[3726] = 8'b00000000;
dat[3727] = 8'b00000000;
dat[3728] = 8'b00000000;
dat[3729] = 8'b00000000;
dat[3730] = 8'b00000000;
dat[3731] = 8'b00000000;
dat[3732] = 8'b00000000;
dat[3733] = 8'b00000000;
dat[3734] = 8'b00000000;
dat[3735] = 8'b00000000;
dat[3736] = 8'b00000000;
dat[3737] = 8'b00000000;
dat[3738] = 8'b00000000;
dat[3739] = 8'b00000000;
dat[3740] = 8'b00000000;
dat[3741] = 8'b00000000;
dat[3742] = 8'b00000000;
dat[3743] = 8'b00000000;
dat[3744] = 8'b00000000;
dat[3745] = 8'b00000000;
dat[3746] = 8'b00000000;
dat[3747] = 8'b00000000;
dat[3748] = 8'b00000000;
dat[3749] = 8'b00000000;
dat[3750] = 8'b00000000;
dat[3751] = 8'b00000000;
dat[3752] = 8'b00000000;
dat[3753] = 8'b00000000;
dat[3754] = 8'b00000000;
dat[3755] = 8'b00000000;
dat[3756] = 8'b00000000;
dat[3757] = 8'b00000000;
dat[3758] = 8'b00000000;
dat[3759] = 8'b00000000;
dat[3760] = 8'b00000000;
dat[3761] = 8'b00000000;
dat[3762] = 8'b00000000;
dat[3763] = 8'b00000000;
dat[3764] = 8'b00000000;
dat[3765] = 8'b00000000;
dat[3766] = 8'b00000000;
dat[3767] = 8'b00000000;
dat[3768] = 8'b00000000;
dat[3769] = 8'b00000000;
dat[3770] = 8'b00000000;
dat[3771] = 8'b00000000;
dat[3772] = 8'b00000000;
dat[3773] = 8'b00000000;
dat[3774] = 8'b00000000;
dat[3775] = 8'b00000000;
dat[3776] = 8'b00000000;
dat[3777] = 8'b00000000;
dat[3778] = 8'b00000000;
dat[3779] = 8'b00000000;
dat[3780] = 8'b00000000;
dat[3781] = 8'b00000000;
dat[3782] = 8'b00000000;
dat[3783] = 8'b00000000;
dat[3784] = 8'b00000000;
dat[3785] = 8'b00000000;
dat[3786] = 8'b00000000;
dat[3787] = 8'b00000000;
dat[3788] = 8'b00000000;
dat[3789] = 8'b00000000;
dat[3790] = 8'b00000000;
dat[3791] = 8'b00000000;
dat[3792] = 8'b00000000;
dat[3793] = 8'b00000000;
dat[3794] = 8'b00000000;
dat[3795] = 8'b00000000;
dat[3796] = 8'b00000000;
dat[3797] = 8'b00000000;
dat[3798] = 8'b00000000;
dat[3799] = 8'b00000000;
dat[3800] = 8'b00000000;
dat[3801] = 8'b00000000;
dat[3802] = 8'b00000000;
dat[3803] = 8'b00000000;
dat[3804] = 8'b00000000;
dat[3805] = 8'b00000000;
dat[3806] = 8'b00000000;
dat[3807] = 8'b00000000;
dat[3808] = 8'b00000000;
dat[3809] = 8'b00000000;
dat[3810] = 8'b00000000;
dat[3811] = 8'b00000000;
dat[3812] = 8'b00000000;
dat[3813] = 8'b00000000;
dat[3814] = 8'b00000000;
dat[3815] = 8'b00000000;
dat[3816] = 8'b00000000;
dat[3817] = 8'b00000000;
dat[3818] = 8'b00000000;
dat[3819] = 8'b00000000;
dat[3820] = 8'b00000000;
dat[3821] = 8'b00000000;
dat[3822] = 8'b00000000;
dat[3823] = 8'b00000000;
dat[3824] = 8'b00000000;
dat[3825] = 8'b00000000;
dat[3826] = 8'b00000000;
dat[3827] = 8'b00000000;
dat[3828] = 8'b00000000;
dat[3829] = 8'b00000000;
dat[3830] = 8'b00000000;
dat[3831] = 8'b00000000;
dat[3832] = 8'b00000000;
dat[3833] = 8'b00000000;
dat[3834] = 8'b00000000;
dat[3835] = 8'b00000000;
dat[3836] = 8'b00000000;
dat[3837] = 8'b00000000;
dat[3838] = 8'b00000000;
dat[3839] = 8'b00000000;
dat[3840] = 8'b00000000;
dat[3841] = 8'b00000000;
dat[3842] = 8'b00000000;
dat[3843] = 8'b00000000;
dat[3844] = 8'b00000000;
dat[3845] = 8'b00000000;
dat[3846] = 8'b00000000;
dat[3847] = 8'b00000000;
dat[3848] = 8'b00000000;
dat[3849] = 8'b00000000;
dat[3850] = 8'b00000000;
dat[3851] = 8'b00000000;
dat[3852] = 8'b00000000;
dat[3853] = 8'b00000000;
dat[3854] = 8'b00000000;
dat[3855] = 8'b00000000;
dat[3856] = 8'b00000000;
dat[3857] = 8'b00000000;
dat[3858] = 8'b00000000;
dat[3859] = 8'b00000000;
dat[3860] = 8'b00000000;
dat[3861] = 8'b00000000;
dat[3862] = 8'b00000000;
dat[3863] = 8'b00000000;
dat[3864] = 8'b00000000;
dat[3865] = 8'b00000000;
dat[3866] = 8'b00000000;
dat[3867] = 8'b00000000;
dat[3868] = 8'b00000000;
dat[3869] = 8'b00000000;
dat[3870] = 8'b00000000;
dat[3871] = 8'b00000000;
dat[3872] = 8'b00000000;
dat[3873] = 8'b00000000;
dat[3874] = 8'b00000000;
dat[3875] = 8'b00000000;
dat[3876] = 8'b00000000;
dat[3877] = 8'b00000000;
dat[3878] = 8'b00000000;
dat[3879] = 8'b00000000;
dat[3880] = 8'b00000000;
dat[3881] = 8'b00000000;
dat[3882] = 8'b00000000;
dat[3883] = 8'b00000000;
dat[3884] = 8'b00000000;
dat[3885] = 8'b00000000;
dat[3886] = 8'b00000000;
dat[3887] = 8'b00000000;
dat[3888] = 8'b00000000;
dat[3889] = 8'b00000000;
dat[3890] = 8'b00000000;
dat[3891] = 8'b00000000;
dat[3892] = 8'b00000000;
dat[3893] = 8'b00000000;
dat[3894] = 8'b00000000;
dat[3895] = 8'b00000000;
dat[3896] = 8'b00000000;
dat[3897] = 8'b00000000;
dat[3898] = 8'b00000000;
dat[3899] = 8'b00000000;
dat[3900] = 8'b00000000;
dat[3901] = 8'b00000000;
dat[3902] = 8'b00000000;
dat[3903] = 8'b00000000;
dat[3904] = 8'b00000000;
dat[3905] = 8'b00000000;
dat[3906] = 8'b00000000;
dat[3907] = 8'b00000000;
dat[3908] = 8'b00000000;
dat[3909] = 8'b00000000;
dat[3910] = 8'b00000000;
dat[3911] = 8'b00000000;
dat[3912] = 8'b00000000;
dat[3913] = 8'b00000000;
dat[3914] = 8'b00000000;
dat[3915] = 8'b00000000;
dat[3916] = 8'b00000000;
dat[3917] = 8'b00000000;
dat[3918] = 8'b00000000;
dat[3919] = 8'b00000000;
dat[3920] = 8'b00000000;
dat[3921] = 8'b00000000;
dat[3922] = 8'b00000000;
dat[3923] = 8'b00000000;
dat[3924] = 8'b00000000;
dat[3925] = 8'b00000000;
dat[3926] = 8'b00000000;
dat[3927] = 8'b00000000;
dat[3928] = 8'b00000000;
dat[3929] = 8'b00000000;
dat[3930] = 8'b00000000;
dat[3931] = 8'b00000000;
dat[3932] = 8'b00000000;
dat[3933] = 8'b00000000;
dat[3934] = 8'b00000000;
dat[3935] = 8'b00000000;
dat[3936] = 8'b00000000;
dat[3937] = 8'b00000000;
dat[3938] = 8'b00000000;
dat[3939] = 8'b00000000;
dat[3940] = 8'b00000000;
dat[3941] = 8'b00000000;
dat[3942] = 8'b00000000;
dat[3943] = 8'b00000000;
dat[3944] = 8'b00000000;
dat[3945] = 8'b00000000;
dat[3946] = 8'b00000000;
dat[3947] = 8'b00000000;
dat[3948] = 8'b00000000;
dat[3949] = 8'b00000000;
dat[3950] = 8'b00000000;
dat[3951] = 8'b00000000;
dat[3952] = 8'b00000000;
dat[3953] = 8'b00000000;
dat[3954] = 8'b00000000;
dat[3955] = 8'b00000000;
dat[3956] = 8'b00000000;
dat[3957] = 8'b00000000;
dat[3958] = 8'b00000000;
dat[3959] = 8'b00000000;
dat[3960] = 8'b00000000;
dat[3961] = 8'b00000000;
dat[3962] = 8'b00000000;
dat[3963] = 8'b00000000;
dat[3964] = 8'b00000000;
dat[3965] = 8'b00000000;
dat[3966] = 8'b00000000;
dat[3967] = 8'b00000000;
dat[3968] = 8'b00000000;
dat[3969] = 8'b00000000;
dat[3970] = 8'b00000000;
dat[3971] = 8'b00000000;
dat[3972] = 8'b00000000;
dat[3973] = 8'b00000000;
dat[3974] = 8'b00000000;
dat[3975] = 8'b00000000;
dat[3976] = 8'b00000000;
dat[3977] = 8'b00000000;
dat[3978] = 8'b00000000;
dat[3979] = 8'b00000000;
dat[3980] = 8'b00000000;
dat[3981] = 8'b00000000;
dat[3982] = 8'b00000000;
dat[3983] = 8'b00000000;
dat[3984] = 8'b00000000;
dat[3985] = 8'b00000000;
dat[3986] = 8'b00000000;
dat[3987] = 8'b00000000;
dat[3988] = 8'b00000000;
dat[3989] = 8'b00000000;
dat[3990] = 8'b00000000;
dat[3991] = 8'b00000000;
dat[3992] = 8'b00000000;
dat[3993] = 8'b00000000;
dat[3994] = 8'b00000000;
dat[3995] = 8'b00000000;
dat[3996] = 8'b00000000;
dat[3997] = 8'b00000000;
dat[3998] = 8'b00000000;
dat[3999] = 8'b00000000;
dat[4000] = 8'b00000000;
dat[4001] = 8'b00000000;
dat[4002] = 8'b00000000;
dat[4003] = 8'b00000000;
dat[4004] = 8'b00000000;
dat[4005] = 8'b00000000;
dat[4006] = 8'b00000000;
dat[4007] = 8'b00000000;
dat[4008] = 8'b00000000;
dat[4009] = 8'b00000000;
dat[4010] = 8'b00000000;
dat[4011] = 8'b00000000;
dat[4012] = 8'b00000000;
dat[4013] = 8'b00000000;
dat[4014] = 8'b00000000;
dat[4015] = 8'b00000000;
dat[4016] = 8'b00000000;
dat[4017] = 8'b00000000;
dat[4018] = 8'b00000000;
dat[4019] = 8'b00000000;
dat[4020] = 8'b00000000;
dat[4021] = 8'b00000000;
dat[4022] = 8'b00000000;
dat[4023] = 8'b00000000;
dat[4024] = 8'b00000000;
dat[4025] = 8'b00000000;
dat[4026] = 8'b00000000;
dat[4027] = 8'b00000000;
dat[4028] = 8'b00000000;
dat[4029] = 8'b00000000;
dat[4030] = 8'b00000000;
dat[4031] = 8'b00000000;
dat[4032] = 8'b00000000;
dat[4033] = 8'b00000000;
dat[4034] = 8'b00000000;
dat[4035] = 8'b00000000;
dat[4036] = 8'b00000000;
dat[4037] = 8'b00000000;
dat[4038] = 8'b00000000;
dat[4039] = 8'b00000000;
dat[4040] = 8'b00000000;
dat[4041] = 8'b00000000;
dat[4042] = 8'b00000000;
dat[4043] = 8'b00000000;
dat[4044] = 8'b00000000;
dat[4045] = 8'b00000000;
dat[4046] = 8'b00000000;
dat[4047] = 8'b00000000;
dat[4048] = 8'b00000000;
dat[4049] = 8'b00000000;
dat[4050] = 8'b00000000;
dat[4051] = 8'b00000000;
dat[4052] = 8'b00000000;
dat[4053] = 8'b00000000;
dat[4054] = 8'b00000000;
dat[4055] = 8'b00000000;
dat[4056] = 8'b00000000;
dat[4057] = 8'b00000000;
dat[4058] = 8'b00000000;
dat[4059] = 8'b00000000;
dat[4060] = 8'b00000000;
dat[4061] = 8'b00000000;
dat[4062] = 8'b00000000;
dat[4063] = 8'b00000000;
dat[4064] = 8'b00000000;
dat[4065] = 8'b00000000;
dat[4066] = 8'b00000000;
dat[4067] = 8'b00000000;
dat[4068] = 8'b00000000;
dat[4069] = 8'b00000000;
dat[4070] = 8'b00000000;
dat[4071] = 8'b00000000;
dat[4072] = 8'b00000000;
dat[4073] = 8'b00000000;
dat[4074] = 8'b00000000;
dat[4075] = 8'b00000000;
dat[4076] = 8'b00000000;
dat[4077] = 8'b00000000;
dat[4078] = 8'b00000000;
dat[4079] = 8'b00000000;
dat[4080] = 8'b00000000;
dat[4081] = 8'b00000000;
dat[4082] = 8'b00000000;
dat[4083] = 8'b00000000;
dat[4084] = 8'b00000000;
dat[4085] = 8'b00000000;
dat[4086] = 8'b00000000;
dat[4087] = 8'b00000000;
dat[4088] = 8'b00000000;
dat[4089] = 8'b00000000;
dat[4090] = 8'b00000000;
dat[4091] = 8'b00000000;
dat[4092] = 8'b00000000;
dat[4093] = 8'b00000000;
dat[4094] = 8'b00000000;
dat[4095] = 8'b00000000;

    end

    // Escreve na memória de dados quando esc_mem é 1
    always @(posedge clock) begin
            if(esc_mem) begin
                dat[dst_mem] <= value[31:24];
                dat[dst_mem + 1] <= value[23:16];
                dat[dst_mem + 2] <= value[15:8];
                dat[dst_mem + 3] <= value[7:0];
            end
    end




    // Atribuições para as saídas
    assign out_dat = {dat[dst_mem], dat[dst_mem + 1], dat[dst_mem + 2], dat[dst_mem + 3]};  // Saída de dados

endmodule
