module MemInst(
    input [31:0] pc,          // endereço de instrução (program counter)
    output [31:0] out_inst,   // saída de instrução (16 bits)
    input clock,
    input stall
);


    // Memória de instruções (256 posições, 8 bits cada)
    reg [7:0] inst [0:8000];

    // Inicialização das memórias

    initial begin //addi,add,sub,jalr e jal(nsalva pc atual, não anterior), sll, or, sra, srl, blt, auipc, lui, lw, sw
    //inst[0] = 32'b00000000-0001_0000-0_000_0001-0_0010011; //addi 2 0 1
    //inst[1] = 32'b0000000_00010_00010_000_00001_0110011; //add 1 0 2
    //inst[2] = 32'b0000000_00001_00000_010_00100_0100011; //sw valor 1 --> 4
    //inst[3] = 32'b000000000100_00000_010_00100_0000011; //lw valor 4 --> 4
    //inst[2] = 32'b00000000000000000010_11111_0010111; //auipc pc + 2
    //inst[2] = 32'b10000000000000000000_11111_0110111; //lui 1 no mais significativo
    //inst[2] = 32'b0000000_00001_00010_100_10100_1100011; //blt pc+10 1 2
    //inst[3] = 32'b0000000_00010_00010_100_10100_1100011; //blt pc+10 1 1
    //inst[2] = 32'b0100000_00010_00001_100_00011_0110011; //sra 3 2 1
    //inst[3] = 32'b0100000_00010_00001_110_00011_0110011; // or 3 2 1
    //inst[4] = 32'b0100000_00010_00001_001_00011_0110011; // sll 3 2 1
    //inst[3] = 32'b0100000_00010_00001_101_00011_0110011; // srl 3 2 1
    //inst[7] = 32'b0100000_00010_00001_011_00011_0110011; //sub 3 2 1
    //inst[3] = 32'b000000001010_00001_000_11111_1100111; //jalr 2 + 10
    //inst[4] = 32'b00000000000000000001_11111_1101111; //jal 1 11111
    //inst[4] = 32'b00000000000000000001_00111_0010111; //aui pc +1, 7
    //inst[5] = 32'b11000000000000000001_11111_0110111; //lui 11...00001 11
/*
// jal test
inst[0] = 8'b00000000;
inst[1] = 8'b00000000;
inst[2] = 8'b00011111;
inst[3] = 8'b11101111;
// addi 2 0 1
inst[4096] = 8'b00000000;
inst[4097] = 8'b00010000;
inst[4098] = 8'b00000001;
inst[4099] = 8'b00010011;
// addi 3 0 2
inst[4100] = 8'b00000000;
inst[4101] = 8'b00100000;
inst[4102] = 8'b00000001;
inst[4103] = 8'b10010011;
// add 1 3 2
inst[4104] = 8'b00000000;
inst[4105] = 8'b00110001;
inst[4106] = 8'b00000000;
inst[4107] = 8'b10110011;
// add 4 3 2
inst[4108] = 8'b00000000;
inst[4109] = 8'b00110001;
inst[4110] = 8'b00000010;
inst[4111] = 8'b00110011;
// add 5 3 2
inst[12] = 8'b00000000;
inst[13] = 8'b00110001;
inst[14] = 8'b00000010;
inst[15] = 8'b10110011;

*/
    //addi 2 0 4
    /*
    inst[0] = 8'b00000000;
    inst[1] = 8'b01000000;
    inst[2] = 8'b00000001;
    inst[3] = 8'b00010011;

    inst[4] = 8'b00000000;
    inst[5] = 8'b00000000;
    inst[6] = 8'b00000000;
    inst[7] = 8'b00000000;

    inst[8] = 8'b00000000;
    inst[9] = 8'b00000000;
    inst[10] = 8'b00000000;
    inst[11] = 8'b00000000;

    inst[12] = 8'b00000000;
    inst[13] = 8'b00000000;
    inst[14] = 8'b00000000;
    inst[15] = 8'b00000000;


    //jalr 2 + 12
    inst[16] = 8'b00000000;
    inst[17] = 8'b1100_0001;
    inst[18] = 8'b0_000_1111;
    inst[19] = 8'b1_1100111;

    inst[20] = 8'b00000000;
    inst[21] = 8'b00000000;
    inst[22] = 8'b00000000;
    inst[23] = 8'b00000000;

    inst[24] = 8'b00000000;
    inst[25] = 8'b00000000;
    inst[26] = 8'b00000000;
    inst[27] = 8'b00000000;

    inst[28] = 8'b00000000;
    inst[29] = 8'b00000000;
    inst[30] = 8'b00000000;
    inst[31] = 8'b00000000;
    */

    // jal test
    /*
inst[0] = 8'b11111000;
inst[1] = 8'b00000000;
inst[2] = 8'b00011111;
inst[3] = 8'b11101111;
// addi 2 0 1
inst[4] = 8'b00000000;
inst[5] = 8'b00010000;
inst[6] = 8'b00000001;
inst[7] = 8'b00010011;
// addi 3 0 2
inst[8] = 8'b00000000;
inst[9] = 8'b00100000;
inst[10] = 8'b00000001;
inst[11] = 8'b10010011;
// add 1 3 2
inst[12] = 8'b00000000;
inst[13] = 8'b00110001;
inst[14] = 8'b00000000;
inst[15] = 8'b10110011;
// add 4 3 2
inst[16] = 8'b00000000;
inst[17] = 8'b00110001;
inst[18] = 8'b00000010;
inst[19] = 8'b00110011;
// add 5 3 2
inst[20] = 8'b00000000;
inst[21] = 8'b00110001;
inst[22] = 8'b00000010;
inst[23] = 8'b10110011;
    */
    /*
    //jal 32 11111
    inst[16] = 8'b00000000;
    inst[17] = 8'b00000010;
    inst[18] = 8'b0000_1111;
    inst[19] = 8'b1_1101111;

    inst[20] = 8'b00000000;
    inst[21] = 8'b00000000;
    inst[22] = 8'b00000000;
    inst[23] = 8'b00000000;

    inst[24] = 8'b00000000;
    inst[25] = 8'b00000000;
    inst[26] = 8'b00000000;
    inst[27] = 8'b00000000;

    inst[28] = 8'b00000000;
    inst[29] = 8'b00000000;
    inst[30] = 8'b00000000;
    inst[31] = 8'b00000000;
    */


    /*
    //addi 2 0 1
    inst[0] = 8'b00000000;
    inst[1] = 8'b00010000;
    inst[2] = 8'b00000001;
    inst[3] = 8'b00010011;

    inst[4] = 8'b00000000;
    inst[5] = 8'b00000000;
    inst[6] = 8'b00000000;
    inst[7] = 8'b00000000;

    inst[8] = 8'b00000000;
    inst[9] = 8'b00000000;
    inst[10] = 8'b00000000;
    inst[11] = 8'b00000000;

    inst[12] = 8'b00000000;
    inst[13] = 8'b00000000;
    inst[14] = 8'b00000000;
    inst[15] = 8'b00000000;

    //add 6 2 1
    inst[16] = 8'b00000000;
    inst[17] = 8'b00010001;
    inst[18] = 8'b00000011;
    inst[19] = 8'b00010011;

    inst[20] = 8'b00000000;
    inst[21] = 8'b00000000;
    inst[22] = 8'b00000000;
    inst[23] = 8'b00000000;

    inst[24] = 8'b00000000;
    inst[25] = 8'b00000000;
    inst[26] = 8'b00000000;
    inst[27] = 8'b00000000;

    inst[28] = 8'b00000000;
    inst[29] = 8'b00000000;
    inst[30] = 8'b00000000;
    inst[31] = 8'b00000000;

    //sub 3 2 1
    inst[32] = 8'b0100000_0;
    inst[33] = 8'b0010_0000;
    inst[34] = 8'b1_011_0001;
    inst[35] = 8'b1_0110011;

    inst[36] = 8'b00000000;
    inst[37] = 8'b00000000;
    inst[38] = 8'b00000000;
    inst[39] = 8'b00000000;

    inst[40] = 8'b00000000;
    inst[41] = 8'b00000000;
    inst[42] = 8'b00000000;
    inst[43] = 8'b00000000;

    inst[44] = 8'b00000000;
    inst[45] = 8'b00000000;
    inst[46] = 8'b00000000;
    inst[47] = 8'b00000000;

    //sw valor 3 --> 4
    inst[48] = 8'b0000000_0;
    inst[49] = 8'b0011_0000;
    inst[50] = 8'b0_010_0010;
    inst[51] = 8'b0_0100011;

    inst[52] = 8'b00000000;
    inst[53] = 8'b00000000;
    inst[54] = 8'b00000000;
    inst[55] = 8'b00000000;

    inst[56] = 8'b00000000;
    inst[57] = 8'b00000000;
    inst[58] = 8'b00000000;
    inst[59] = 8'b00000000;

    inst[60] = 8'b00000000;
    inst[61] = 8'b00000000;
    inst[62] = 8'b00000000;
    inst[63] = 8'b00000000;

    //lw valor 4 --> 4
    inst[64] = 8'b00000000;
    inst[65] = 8'b0100_0000;
    inst[66] = 8'b0_010_0010;
    inst[67] = 8'b0_0000011;

    inst[68] = 8'b00000000;
    inst[69] = 8'b00000000;
    inst[70] = 8'b00000000;
    inst[71] = 8'b00000000;

    inst[72] = 8'b00000000;
    inst[73] = 8'b00000000;
    inst[74] = 8'b00000000;
    inst[75] = 8'b00000000;

    inst[76] = 8'b00000000;
    inst[77] = 8'b00000000;
    inst[78] = 8'b00000000;
    inst[79] = 8'b00000000;

    //auipc pc + 2 --> 31
    inst[80] = 8'b00000000;
    inst[81] = 8'b00000000;
    inst[82] = 8'b0010_1111;
    inst[83] = 8'b1_0010111;

    inst[84] = 8'b00000000;
    inst[85] = 8'b00000000;
    inst[86] = 8'b00000000;
    inst[87] = 8'b00000000;

    inst[88] = 8'b00000000;
    inst[89] = 8'b00000000;
    inst[90] = 8'b00000000;
    inst[91] = 8'b00000000;

    inst[92] = 8'b00000000;
    inst[93] = 8'b00000000;
    inst[94] = 8'b00000000;
    inst[95] = 8'b00000000;

    //lui 1 no mais significativo
    inst[96] = 8'b10000000;
    inst[97] = 8'b00000000;
    inst[98] = 8'b0000_1111;
    inst[99] = 8'b1_0110111;

    inst[100] = 8'b00000000;
    inst[101] = 8'b00000000;
    inst[102] = 8'b00000000;
    inst[103] = 8'b00000000;

    inst[104] = 8'b00000000;
    inst[105] = 8'b00000000;
    inst[106] = 8'b00000000;
    inst[107] = 8'b00000000;

    inst[108] = 8'b00000000;
    inst[109] = 8'b00000000;
    inst[110] = 8'b00000000;
    inst[111] = 8'b00000000;

    //blt pc+10 1 2
    inst[112] = 8'b0000000_0;
    inst[113] = 8'b0001_0001;
    inst[114] = 8'b0_100_1000;
    inst[115] = 8'b0_1100011;

    inst[116] = 8'b00000000;
    inst[117] = 8'b00000000;
    inst[118] = 8'b00000000;
    inst[119] = 8'b00000000;

    inst[120] = 8'b00000000;
    inst[121] = 8'b00000000;
    inst[122] = 8'b00000000;
    inst[123] = 8'b00000000;

    inst[124] = 8'b00000000;
    inst[125] = 8'b00000000;
    inst[126] = 8'b00000000;
    inst[127] = 8'b00000000;

    //blt pc+10 1 1
    inst[128] = 8'b0000000_0;
    inst[129] = 8'b001_00000_;
    inst[130] = 8'b010_01000;
    inst[131] = 8'b0_1100011;

    inst[132] = 8'b00000000;
    inst[133] = 8'b00000000;
    inst[134] = 8'b00000000;
    inst[135]= 8'b00000000;

    inst[136] = 8'b00000000;
    inst[137] = 8'b00000000;
    inst[138] = 8'b00000000;
    inst[139] = 8'b00000000;

    inst[140] = 8'b00000000;
    inst[141] = 8'b00000000;
    inst[142] = 8'b00000000;
    inst[143] = 8'b00000000;
    */
        // ... (inicialize o restante das posições com 0)

        // Instruções já fornecidas
inst[0] = 8'b11111110;
inst[1] = 8'b00000001;
inst[2] = 8'b00000001;
inst[3] = 8'b00010011;

inst[4] = 8'b0000000_0;
inst[5] = 8'b0001_0001;
inst[6] = 8'b0_010_1110;
inst[7] = 8'b0_0100011;

inst[8] = 8'b00000000;
inst[9] = 8'b10000001;
inst[10] = 8'b00101100;
inst[11] = 8'b00100011;
inst[12] = 8'b00000010;
inst[13] = 8'b00000001;
inst[14] = 8'b00000100;
inst[15] = 8'b00010011;
inst[16] = 8'b00000000;
inst[17] = 8'b00000000;
inst[18] = 8'b00000111;
inst[19] = 8'b10110111;
inst[20] = 8'b00000000;
inst[21] = 8'b00000111;
inst[22] = 8'b10000111;
inst[23] = 8'b10010011;
inst[24] = 8'b00000000;
inst[25] = 8'b00000111;
inst[26] = 8'b10100110;
inst[27] = 8'b00000011;
inst[28] = 8'b00000000;
inst[29] = 8'b01000111;
inst[30] = 8'b10100110;
inst[31] = 8'b10000011;
inst[32] = 8'b00000000;
inst[33] = 8'b10000111;
inst[34] = 8'b10100111;
inst[35] = 8'b00000011;
inst[36] = 8'b00000000;
inst[37] = 8'b11000111;
inst[38] = 8'b10100111;
inst[39] = 8'b10000011;
inst[40] = 8'b11111110;
inst[41] = 8'b11000100;
inst[42] = 8'b00100000;
inst[43] = 8'b00100011;
inst[44] = 8'b11111110;
inst[45] = 8'b11010100;
inst[46] = 8'b00100010;
inst[47] = 8'b00100011;
inst[48] = 8'b11111110;
inst[49] = 8'b11100100;
inst[50] = 8'b00100100;
inst[51] = 8'b00100011;
inst[52] = 8'b11111110;
inst[53] = 8'b11110100;
inst[54] = 8'b00100110;
inst[55] = 8'b00100011;
inst[56] = 8'b11111110;
inst[57] = 8'b00000100;
inst[58] = 8'b00000111;
inst[59] = 8'b10010011;
inst[60] = 8'b00000000;
inst[61] = 8'b00110000;
inst[62] = 8'b00000110;
inst[63] = 8'b00010011;
inst[64] = 8'b00000000;
inst[65] = 8'b00000000;
inst[66] = 8'b00000101;
inst[67] = 8'b10010011;
inst[68] = 8'b00000000;
inst[69] = 8'b00000111;
inst[70] = 8'b10000101;
inst[71] = 8'b00010011;
inst[72] = 8'b00000000;
inst[73] = 8'b00000000;
inst[74] = 8'b00000000;
inst[75] = 8'b10010111;

inst[76] = 8'b00111000;
inst[77] = 8'b1100_0000;
inst[78] = 8'b1_000_0000;
inst[79] = 8'b1_1100111;

inst[80] = 8'b00000000;
inst[81] = 8'b00000000;
inst[82] = 8'b00000111;
inst[83] = 8'b10010011;
inst[84] = 8'b00000000;
inst[85] = 8'b00000111;
inst[86] = 8'b10000101;
inst[87] = 8'b00010011;
inst[88] = 8'b00000001;
inst[89] = 8'b11000001;
inst[90] = 8'b00100000;
inst[91] = 8'b10000011;
inst[92] = 8'b00000001;
inst[93] = 8'b10000001;
inst[94] = 8'b00100100;
inst[95] = 8'b00000011;
inst[96] = 8'b00000010;
inst[97] = 8'b00000001;
inst[98] = 8'b00000001;
inst[99] = 8'b00010011;

inst[100] = 8'b01111111;
inst[101] = 8'b11111111;
inst[102] = 8'b1111_0000;
inst[103] = 8'b0_1100111;

inst[104] = 8'b11111010;
inst[105] = 8'b00000001;
inst[106] = 8'b00000001;
inst[107] = 8'b00010011;
inst[108] = 8'b00000100;
inst[109] = 8'b10000001;
inst[110] = 8'b00101110;
inst[111] = 8'b00100011;
inst[112] = 8'b00000101;
inst[113] = 8'b00100001;
inst[114] = 8'b00101100;
inst[115] = 8'b00100011;
inst[116] = 8'b00000101;
inst[117] = 8'b00110001;
inst[118] = 8'b00101010;
inst[119] = 8'b00100011;
inst[120] = 8'b00000101;
inst[121] = 8'b01000001;
inst[122] = 8'b00101000;
inst[123] = 8'b00100011;
inst[124] = 8'b00000101;
inst[125] = 8'b01010001;
inst[126] = 8'b00100110;
inst[127] = 8'b00100011;
inst[128] = 8'b00000101;
inst[129] = 8'b01100001;
inst[130] = 8'b00100100;
inst[131] = 8'b00100011;
inst[132] = 8'b00000101;
inst[133] = 8'b01110001;
inst[134] = 8'b00100010;
inst[135] = 8'b00100011;
inst[136] = 8'b00000110;
inst[137] = 8'b00000001;
inst[138] = 8'b00000100;
inst[139] = 8'b00010011;
inst[140] = 8'b11111010;
inst[141] = 8'b10100100;
inst[142] = 8'b00100110;
inst[143] = 8'b00100011;
inst[144] = 8'b11111010;
inst[145] = 8'b10110100;
inst[146] = 8'b00100100;
inst[147] = 8'b00100011;
inst[148] = 8'b11111010;
inst[149] = 8'b11000100;
inst[150] = 8'b00100010;
inst[151] = 8'b00100011;
inst[152] = 8'b11111010;
inst[153] = 8'b11010100;
inst[154] = 8'b00100000;
inst[155] = 8'b00100011;
inst[156] = 8'b00000000;
inst[157] = 8'b00000001;
inst[158] = 8'b00000110;
inst[159] = 8'b10010011;
inst[160] = 8'b00000000;
inst[161] = 8'b00000110;
inst[162] = 8'b10000101;
inst[163] = 8'b10010011;
inst[164] = 8'b11111010;
inst[165] = 8'b01000100;
inst[166] = 8'b00100110;
inst[167] = 8'b00000011;
inst[168] = 8'b11111010;
inst[169] = 8'b10000100;
inst[170] = 8'b00100110;
inst[171] = 8'b10000011;
//
inst[172] = 8'b01000000;
inst[173] = 8'b11010110;
inst[174] = 8'b11000110;
inst[175] = 8'b10110011;
inst[176] = 8'b00000000;
inst[177] = 8'b00010110;
inst[178] = 8'b10000110;
inst[179] = 8'b10010011;
inst[180] = 8'b11111100;
inst[181] = 8'b11010100;
inst[182] = 8'b00101000;
inst[183] = 8'b00100011;
inst[184] = 8'b11111010;
inst[185] = 8'b00000100;
inst[186] = 8'b00100110;
inst[187] = 8'b00000011;
inst[188] = 8'b11111010;
inst[189] = 8'b01000100;
inst[190] = 8'b00100110;
inst[191] = 8'b10000011;
//
inst[192] = 8'b01000000;
inst[193] = 8'b11010110;
inst[194] = 8'b00110110;
inst[195] = 8'b10110011;
inst[196] = 8'b11111100;
inst[197] = 8'b11010100;
inst[198] = 8'b00100110;
inst[199] = 8'b00100011;
inst[200] = 8'b11111101;
inst[201] = 8'b00000100;
inst[202] = 8'b00100110;
inst[203] = 8'b10000011;
inst[204] = 8'b11111111;
inst[205] = 8'b11110110;
inst[206] = 8'b10000110;
inst[207] = 8'b00010011;
inst[208] = 8'b11111100;
inst[209] = 8'b11000100;
inst[210] = 8'b00100100;
inst[211] = 8'b00100011;
inst[212] = 8'b00000000;
inst[213] = 8'b00000110;
inst[214] = 8'b10000110;
inst[215] = 8'b00010011;
inst[216] = 8'b00000000;
inst[217] = 8'b00000110;
inst[218] = 8'b00001011;
inst[219] = 8'b00010011;
inst[220] = 8'b00000000;
inst[221] = 8'b00000000;
inst[222] = 8'b00001011;
inst[223] = 8'b10010011;
inst[224] = 8'b00000001;
inst[225] = 8'b10111011;
inst[226] = 8'b01010110;
inst[227] = 8'b00010011;
inst[228] = 8'b00000000;
inst[229] = 8'b01011011;
inst[230] = 8'b10011110;
inst[231] = 8'b10010011;
inst[232] = 8'b00000001;
inst[233] = 8'b11010110;
inst[234] = 8'b01101110;
inst[235] = 8'b10110011;
inst[236] = 8'b00000000;
inst[237] = 8'b01011011;
inst[238] = 8'b00011110;
inst[239] = 8'b00010011;
inst[240] = 8'b00000000;
inst[241] = 8'b00000110;
inst[242] = 8'b10000110;
inst[243] = 8'b00010011;
inst[244] = 8'b00000000;
inst[245] = 8'b00000110;
inst[246] = 8'b00001010;
inst[247] = 8'b00010011;
inst[248] = 8'b00000000;
inst[249] = 8'b00000000;
inst[250] = 8'b00001010;
inst[251] = 8'b10010011;
inst[252] = 8'b00000001;
inst[253] = 8'b10111010;
inst[254] = 8'b01010110;
inst[255] = 8'b00010011;
inst[256] = 8'b00000000;
inst[257] = 8'b01011010;
inst[258] = 8'b10010011;
inst[259] = 8'b10010011;
inst[260] = 8'b00000000;
inst[261] = 8'b01110110;
inst[262] = 8'b01100011;
inst[263] = 8'b10110011;
inst[264] = 8'b00000000;
inst[265] = 8'b01011010;
inst[266] = 8'b00010011;
inst[267] = 8'b00010011;
inst[268] = 8'b00000000;
inst[269] = 8'b00100110;
inst[270] = 8'b10010110;
inst[271] = 8'b10010011;
inst[272] = 8'b00000000;
inst[273] = 8'b11110110;
inst[274] = 8'b10000110;
inst[275] = 8'b10010011;
inst[276] = 8'b00000000;
inst[277] = 8'b01000110;
inst[278] = 8'b11010110;
inst[279] = 8'b10010011;
inst[280] = 8'b00000000;
inst[281] = 8'b01000110;
inst[282] = 8'b10010110;
inst[283] = 8'b10010011;
//
inst[284] = 8'b01000000;
inst[285] = 8'b11010001;
inst[286] = 8'b00110001;
inst[287] = 8'b00110011;
inst[288] = 8'b00000000;
inst[289] = 8'b00000001;
inst[290] = 8'b00000110;
inst[291] = 8'b10010011;
inst[292] = 8'b00000000;
inst[293] = 8'b00110110;
inst[294] = 8'b10000110;
inst[295] = 8'b10010011;
inst[296] = 8'b00000000;
inst[297] = 8'b00100110;
inst[298] = 8'b11010110;
inst[299] = 8'b10010011;
inst[300] = 8'b00000000;
inst[301] = 8'b00100110;
inst[302] = 8'b10010110;
inst[303] = 8'b10010011;
inst[304] = 8'b11111100;
inst[305] = 8'b11010100;
inst[306] = 8'b00100010;
inst[307] = 8'b00100011;
inst[308] = 8'b11111100;
inst[309] = 8'b11000100;
inst[310] = 8'b00100110;
inst[311] = 8'b10000011;
inst[312] = 8'b11111111;
inst[313] = 8'b11110110;
inst[314] = 8'b10000110;
inst[315] = 8'b00010011;
inst[316] = 8'b11111100;
inst[317] = 8'b11000100;
inst[318] = 8'b00100000;
inst[319] = 8'b00100011;
inst[320] = 8'b00000000;
inst[321] = 8'b00000110;
inst[322] = 8'b10000110;
inst[323] = 8'b00010011;
inst[324] = 8'b00000000;
inst[325] = 8'b00000110;
inst[326] = 8'b00001001;
inst[327] = 8'b00010011;
inst[328] = 8'b00000000;
inst[329] = 8'b00000000;
inst[330] = 8'b00001001;
inst[331] = 8'b10010011;
inst[332] = 8'b00000001;
inst[333] = 8'b10111001;
inst[334] = 8'b01010110;
inst[335] = 8'b00010011;
inst[336] = 8'b00000000;
inst[337] = 8'b01011001;
inst[338] = 8'b10011000;
inst[339] = 8'b10010011;
inst[340] = 8'b00000001;
inst[341] = 8'b00010110;
inst[342] = 8'b01101000;
inst[343] = 8'b10110011;
inst[344] = 8'b00000000;
inst[345] = 8'b01011001;
inst[346] = 8'b00011000;
inst[347] = 8'b00010011;
inst[348] = 8'b00000000;
inst[349] = 8'b00000110;
inst[350] = 8'b10000110;
inst[351] = 8'b00010011;
inst[352] = 8'b00000000;
inst[353] = 8'b00000110;
inst[354] = 8'b00001111;
inst[355] = 8'b00010011;
inst[356] = 8'b00000000;
inst[357] = 8'b00000000;
inst[358] = 8'b00001111;
inst[359] = 8'b10010011;
inst[360] = 8'b00000001;
inst[361] = 8'b10111111;
inst[362] = 8'b01010110;
inst[363] = 8'b00010011;
inst[364] = 8'b00000000;
inst[365] = 8'b01011111;
inst[366] = 8'b10010111;
inst[367] = 8'b10010011;
inst[368] = 8'b00000000;
inst[369] = 8'b11110110;
inst[370] = 8'b01100111;
inst[371] = 8'b10110011;
inst[372] = 8'b00000000;
inst[373] = 8'b01011111;
inst[374] = 8'b00010111;
inst[375] = 8'b00010011;
inst[376] = 8'b00000000;
inst[377] = 8'b00000110;
inst[378] = 8'b10000111;
inst[379] = 8'b10010011;
inst[380] = 8'b00000000;
inst[381] = 8'b00100111;
inst[382] = 8'b10010111;
inst[383] = 8'b10010011;
inst[384] = 8'b00000000;
inst[385] = 8'b11110111;
inst[386] = 8'b10000111;
inst[387] = 8'b10010011;
inst[388] = 8'b00000000;
inst[389] = 8'b01000111;
inst[390] = 8'b11010111;
inst[391] = 8'b10010011;
inst[392] = 8'b00000000;
inst[393] = 8'b01000111;
inst[394] = 8'b10010111;
inst[395] = 8'b10010011;
//
inst[396] = 8'b01000000;
inst[397] = 8'b11110001;
inst[398] = 8'b00110001;
inst[399] = 8'b00110011;
inst[400] = 8'b00000000;
inst[401] = 8'b00000001;
inst[402] = 8'b00000111;
inst[403] = 8'b10010011;
inst[404] = 8'b00000000;
inst[405] = 8'b00110111;
inst[406] = 8'b10000111;
inst[407] = 8'b10010011;
inst[408] = 8'b00000000;
inst[409] = 8'b00100111;
inst[410] = 8'b11010111;
inst[411] = 8'b10010011;
inst[412] = 8'b00000000;
inst[413] = 8'b00100111;
inst[414] = 8'b10010111;
inst[415] = 8'b10010011;
inst[416] = 8'b11111010;
inst[417] = 8'b11110100;
inst[418] = 8'b00101110;
inst[419] = 8'b00100011;
inst[420] = 8'b11111100;
inst[421] = 8'b00000100;
inst[422] = 8'b00101010;
inst[423] = 8'b00100011;
inst[424] = 8'b00000100;
inst[425] = 8'b00000000;
inst[426] = 8'b00000000;
inst[427] = 8'b01101111;
inst[428] = 8'b11111010;
inst[429] = 8'b10000100;
inst[430] = 8'b00100111;
inst[431] = 8'b00000011;
inst[432] = 8'b11111101;
inst[433] = 8'b01000100;
inst[434] = 8'b00100111;
inst[435] = 8'b10000011;

inst[436] = 8'b00000000;
inst[437] = 8'b11110111;
inst[438] = 8'b00000111;
inst[439] = 8'b1_0110011;

inst[440] = 8'b00000000;
inst[441] = 8'b0010_0111;
inst[442] = 8'b1_001_0111;
inst[443] = 8'b1_0010011;

inst[444] = 8'b11111010;
inst[445] = 8'b11000100;
inst[446] = 8'b00100111;
inst[447] = 8'b00000011;
inst[448] = 8'b00000000;
inst[449] = 8'b11110111;
inst[450] = 8'b00000111;
inst[451] = 8'b10110011;
inst[452] = 8'b00000000;
inst[453] = 8'b00000111;
inst[454] = 8'b10100111;
inst[455] = 8'b00000011;
inst[456] = 8'b11111100;
inst[457] = 8'b01000100;
inst[458] = 8'b00100110;
inst[459] = 8'b10000011;
inst[460] = 8'b11111101;
inst[461] = 8'b01000100;
inst[462] = 8'b00100111;
inst[463] = 8'b10000011;
inst[464] = 8'b00000000;
inst[465] = 8'b00100111;
inst[466] = 8'b10010111;
inst[467] = 8'b10010011;
inst[468] = 8'b00000000;
inst[469] = 8'b11110110;
inst[470] = 8'b10000111;
inst[471] = 8'b10110011;
inst[472] = 8'b00000000;
inst[473] = 8'b11100111;
inst[474] = 8'b10100000;
inst[475] = 8'b00100011;
inst[476] = 8'b11111101;
inst[477] = 8'b01000100;
inst[478] = 8'b00100111;
inst[479] = 8'b10000011;
inst[480] = 8'b00000000;
inst[481] = 8'b00010111;
inst[482] = 8'b10000111;
inst[483] = 8'b10010011;
inst[484] = 8'b11111100;
inst[485] = 8'b11110100;
inst[486] = 8'b00101010;
inst[487] = 8'b00100011;
inst[488] = 8'b11111101;
inst[489] = 8'b01000100;
inst[490] = 8'b00100111;
inst[491] = 8'b00000011;
inst[492] = 8'b11111101;
inst[493] = 8'b00000100;
inst[494] = 8'b00100111;
inst[495] = 8'b10000011;
inst[496] = 8'b11111010;
inst[497] = 8'b11110111;
inst[498] = 8'b01001110;
inst[499] = 8'b11100011;
inst[500] = 8'b11111100;
inst[501] = 8'b00000100;
inst[502] = 8'b00101100;
inst[503] = 8'b00100011;
inst[504] = 8'b00000100;
inst[505] = 8'b01000000;
inst[506] = 8'b00000000;
inst[507] = 8'b01101111;
inst[508] = 8'b11111010;
inst[509] = 8'b01000100;
inst[510] = 8'b00100111;
inst[511] = 8'b10000011;
inst[512] = 8'b00000000;
inst[513] = 8'b00010111;
inst[514] = 8'b10000111;
inst[515] = 8'b00010011;
inst[516] = 8'b11111101;
inst[517] = 8'b10000100;
inst[518] = 8'b00100111;
inst[519] = 8'b10000011;
inst[520] = 8'b00000000;
inst[521] = 8'b11110111;
inst[522] = 8'b00000111;
inst[523] = 8'b10110011;
inst[524] = 8'b00000000;
inst[525] = 8'b00100111;
inst[526] = 8'b10010111;
inst[527] = 8'b10010011;
inst[528] = 8'b11111010;
inst[529] = 8'b11000100;
inst[530] = 8'b00100111;
inst[531] = 8'b00000011;
inst[532] = 8'b00000000;
inst[533] = 8'b11110111;
inst[534] = 8'b00000111;
inst[535] = 8'b10110011;
inst[536] = 8'b00000000;
inst[537] = 8'b00000111;
inst[538] = 8'b10100111;
inst[539] = 8'b00000011;
inst[540] = 8'b11111011;
inst[541] = 8'b11000100;
inst[542] = 8'b00100110;
inst[543] = 8'b10000011;
inst[544] = 8'b11111101;
inst[545] = 8'b10000100;
inst[546] = 8'b00100111;
inst[547] = 8'b10000011;
inst[548] = 8'b00000000;
inst[549] = 8'b00100111;
inst[550] = 8'b10010111;
inst[551] = 8'b10010011;
inst[552] = 8'b00000000;
inst[553] = 8'b11110110;
inst[554] = 8'b10000111;
inst[555] = 8'b10110011;
inst[556] = 8'b00000000;
inst[557] = 8'b11100111;
inst[558] = 8'b10100000;
inst[559] = 8'b00100011;
inst[560] = 8'b11111101;
inst[561] = 8'b10000100;
inst[562] = 8'b00100111;
inst[563] = 8'b10000011;
inst[564] = 8'b00000000;
inst[565] = 8'b00010111;
inst[566] = 8'b10000111;
inst[567] = 8'b10010011;
inst[568] = 8'b11111100;
inst[569] = 8'b11110100;
inst[570] = 8'b00101100;
inst[571] = 8'b00100011;
inst[572] = 8'b11111101;
inst[573] = 8'b10000100;
inst[574] = 8'b00100111;
inst[575] = 8'b00000011;
inst[576] = 8'b11111100;
inst[577] = 8'b11000100;
inst[578] = 8'b00100111;
inst[579] = 8'b10000011;
inst[580] = 8'b11111010;
inst[581] = 8'b11110111;
inst[582] = 8'b01001100;
inst[583] = 8'b11100011;
inst[584] = 8'b11111100;
inst[585] = 8'b00000100;
inst[586] = 8'b00101010;
inst[587] = 8'b00100011;
inst[588] = 8'b11111100;
inst[589] = 8'b00000100;
inst[590] = 8'b00101100;
inst[591] = 8'b00100011;
inst[592] = 8'b11111010;
inst[593] = 8'b10000100;
inst[594] = 8'b00100111;
inst[595] = 8'b10000011;
inst[596] = 8'b11111100;
inst[597] = 8'b11110100;
inst[598] = 8'b00101110;
inst[599] = 8'b00100011;
inst[600] = 8'b00001010;
inst[601] = 8'b01000000;
inst[602] = 8'b00000000;
inst[603] = 8'b01101111;
inst[604] = 8'b11111100;
inst[605] = 8'b01000100;
inst[606] = 8'b00100111;
inst[607] = 8'b00000011;
inst[608] = 8'b11111101;
inst[609] = 8'b01000100;
inst[610] = 8'b00100111;
inst[611] = 8'b10000011;
inst[612] = 8'b00000000;
inst[613] = 8'b00100111;
inst[614] = 8'b10010111;
inst[615] = 8'b10010011;
inst[616] = 8'b00000000;
inst[617] = 8'b11110111;
inst[618] = 8'b00000111;
inst[619] = 8'b10110011;
inst[620] = 8'b00000000;
inst[621] = 8'b00000111;
inst[622] = 8'b10100111;
inst[623] = 8'b00000011;
inst[624] = 8'b11111011;
inst[625] = 8'b11000100;
inst[626] = 8'b00100110;
inst[627] = 8'b10000011;
inst[628] = 8'b11111101;
inst[629] = 8'b10000100;
inst[630] = 8'b00100111;
inst[631] = 8'b10000011;
inst[632] = 8'b00000000;
inst[633] = 8'b00100111;
inst[634] = 8'b10010111;
inst[635] = 8'b10010011;
inst[636] = 8'b00000000;
inst[637] = 8'b11110110;
inst[638] = 8'b10000111;
inst[639] = 8'b10110011;
inst[640] = 8'b00000000;
inst[641] = 8'b00000111;
inst[642] = 8'b10100111;
inst[643] = 8'b10000011;
inst[644] = 8'b00000100;
inst[645] = 8'b11100111;
inst[646] = 8'b11000000;
inst[647] = 8'b01100011;
inst[648] = 8'b11111101;
inst[649] = 8'b01000100;
inst[650] = 8'b00100111;
inst[651] = 8'b10000011;
inst[652] = 8'b00000000;
inst[653] = 8'b00010111;
inst[654] = 8'b10000111;
inst[655] = 8'b00010011;
inst[656] = 8'b11111100;
inst[657] = 8'b11100100;
inst[658] = 8'b00101010;
inst[659] = 8'b00100011;
inst[660] = 8'b11111101;
inst[661] = 8'b11000100;
inst[662] = 8'b00100111;
inst[663] = 8'b00000011;
inst[664] = 8'b00000000;
inst[665] = 8'b00010111;
inst[666] = 8'b00000110;
inst[667] = 8'b10010011;
inst[668] = 8'b11111100;
inst[669] = 8'b11010100;
inst[670] = 8'b00101110;
inst[671] = 8'b00100011;
inst[672] = 8'b00000000;
inst[673] = 8'b00100111;
inst[674] = 8'b00010111;
inst[675] = 8'b00010011;
inst[676] = 8'b11111010;
inst[677] = 8'b11000100;
inst[678] = 8'b00100110;
inst[679] = 8'b10000011;
inst[680] = 8'b00000000;
inst[681] = 8'b11100110;
inst[682] = 8'b10000111;
inst[683] = 8'b00110011;
inst[684] = 8'b11111100;
inst[685] = 8'b01000100;
inst[686] = 8'b00100110;
inst[687] = 8'b10000011;
inst[688] = 8'b00000000;
inst[689] = 8'b00100111;
inst[690] = 8'b10010111;
inst[691] = 8'b10010011;
inst[692] = 8'b00000000;
inst[693] = 8'b11110110;
inst[694] = 8'b10000111;
inst[695] = 8'b10110011;
inst[696] = 8'b00000000;
inst[697] = 8'b00000111;
inst[698] = 8'b10100111;
inst[699] = 8'b10000011;
inst[700] = 8'b00000000;
inst[701] = 8'b11110111;
inst[702] = 8'b00100000;
inst[703] = 8'b00100011;
inst[704] = 8'b00000011;
inst[705] = 8'b11000000;
inst[706] = 8'b00000000;
inst[707] = 8'b01101111;
inst[708] = 8'b11111101;
inst[709] = 8'b10000100;
inst[710] = 8'b00100111;
inst[711] = 8'b10000011;
inst[712] = 8'b00000000;
inst[713] = 8'b00010111;
inst[714] = 8'b10000111;
inst[715] = 8'b00010011;
inst[716] = 8'b11111100;
inst[717] = 8'b11100100;
inst[718] = 8'b00101100;
inst[719] = 8'b00100011;
inst[720] = 8'b11111101;
inst[721] = 8'b11000100;
inst[722] = 8'b00100111;
inst[723] = 8'b00000011;
inst[724] = 8'b00000000;
inst[725] = 8'b00010111;
inst[726] = 8'b00000110;
inst[727] = 8'b10010011;
inst[728] = 8'b11111100;
inst[729] = 8'b11010100;
inst[730] = 8'b00101110;
inst[731] = 8'b00100011;
inst[732] = 8'b00000000;
inst[733] = 8'b00100111;
inst[734] = 8'b00010111;
inst[735] = 8'b00010011;
inst[736] = 8'b11111010;
inst[737] = 8'b11000100;
inst[738] = 8'b00100110;
inst[739] = 8'b10000011;
inst[740] = 8'b00000000;
inst[741] = 8'b11100110;
inst[742] = 8'b10000111;
inst[743] = 8'b00110011;
inst[744] = 8'b11111011;
inst[745] = 8'b11000100;
inst[746] = 8'b00100110;
inst[747] = 8'b10000011;
inst[748] = 8'b00000000;
inst[749] = 8'b00100111;
inst[750] = 8'b10010111;
inst[751] = 8'b10010011;
inst[752] = 8'b00000000;
inst[753] = 8'b11110110;
inst[754] = 8'b10000111;
inst[755] = 8'b10110011;
inst[756] = 8'b00000000;
inst[757] = 8'b00000111;
inst[758] = 8'b10100111;
inst[759] = 8'b10000011;
inst[760] = 8'b00000000;
inst[761] = 8'b11110111;
inst[762] = 8'b00100000;
inst[763] = 8'b00100011;
inst[764] = 8'b11111101;
inst[765] = 8'b01000100;
inst[766] = 8'b00100111;
inst[767] = 8'b00000011;
inst[768] = 8'b11111101;
inst[769] = 8'b00000100;
inst[770] = 8'b00100111;
inst[771] = 8'b10000011;
// 0000010_01111_01110_101_01100_1100011
inst[772] = 8'b00000100;
inst[773] = 8'b11100111;
inst[774] = 8'b11000110;
inst[775] = 8'b01100011;
inst[776] = 8'b11111101;
inst[777] = 8'b10000100;
inst[778] = 8'b00100111;
inst[779] = 8'b00000011;
inst[780] = 8'b11111100;
inst[781] = 8'b11000100;
inst[782] = 8'b00100111;
inst[783] = 8'b10000011;
inst[784] = 8'b11110100;
inst[785] = 8'b11110111;
inst[786] = 8'b01000110;
inst[787] = 8'b11100011;
inst[788] = 8'b00000011;
inst[789] = 8'b11000000;
inst[790] = 8'b00000000;
inst[791] = 8'b01101111;
inst[792] = 8'b11111101;
inst[793] = 8'b01000100;
inst[794] = 8'b00100111;
inst[795] = 8'b10000011;
inst[796] = 8'b00000000;
inst[797] = 8'b00010111;
inst[798] = 8'b10000111;
inst[799] = 8'b00010011;
inst[800] = 8'b11111100;
inst[801] = 8'b11100100;
inst[802] = 8'b00101010;
inst[803] = 8'b00100011;
inst[804] = 8'b11111101;
inst[805] = 8'b11000100;
inst[806] = 8'b00100111;
inst[807] = 8'b00000011;
inst[808] = 8'b00000000;
inst[809] = 8'b00010111;
inst[810] = 8'b00000110;
inst[811] = 8'b10010011;
inst[812] = 8'b11111100;
inst[813] = 8'b11010100;
inst[814] = 8'b00101110;
inst[815] = 8'b00100011;
inst[816] = 8'b00000000;
inst[817] = 8'b00100111;
inst[818] = 8'b00010111;
inst[819] = 8'b00010011;
inst[820] = 8'b11111010;
inst[821] = 8'b11000100;
inst[822] = 8'b00100110;
inst[823] = 8'b10000011;
inst[824] = 8'b00000000;
inst[825] = 8'b11100110;
inst[826] = 8'b10000111;
inst[827] = 8'b00110011;
inst[828] = 8'b11111100;
inst[829] = 8'b01000100;
inst[830] = 8'b00100110;
inst[831] = 8'b10000011;
inst[832] = 8'b00000000;
inst[833] = 8'b00100111;
inst[834] = 8'b10010111;
inst[835] = 8'b10010011;
inst[836] = 8'b00000000;
inst[837] = 8'b11110110;
inst[838] = 8'b10000111;
inst[839] = 8'b10110011;
inst[840] = 8'b00000000;
inst[841] = 8'b00000111;
inst[842] = 8'b10100111;
inst[843] = 8'b10000011;
inst[844] = 8'b00000000;
inst[845] = 8'b11110111;
inst[846] = 8'b00100000;
inst[847] = 8'b00100011;
inst[848] = 8'b11111101;
inst[849] = 8'b01000100;
inst[850] = 8'b00100111;
inst[851] = 8'b00000011;
inst[852] = 8'b11111101;
inst[853] = 8'b00000100;
inst[854] = 8'b00100111;
inst[855] = 8'b10000011;
inst[856] = 8'b11111100;
inst[857] = 8'b11110111;
inst[858] = 8'b01000000;
inst[859] = 8'b11100011;
inst[860] = 8'b00000011;
inst[861] = 8'b11000000;
inst[862] = 8'b00000000;
inst[863] = 8'b01101111;
inst[864] = 8'b11111101;
inst[865] = 8'b10000100;
inst[866] = 8'b00100111;
inst[867] = 8'b10000011;
inst[868] = 8'b00000000;
inst[869] = 8'b00010111;
inst[870] = 8'b10000111;
inst[871] = 8'b00010011;
inst[872] = 8'b11111100;
inst[873] = 8'b11100100;
inst[874] = 8'b00101100;
inst[875] = 8'b00100011;
inst[876] = 8'b11111101;
inst[877] = 8'b11000100;
inst[878] = 8'b00100111;
inst[879] = 8'b00000011;
inst[880] = 8'b00000000;
inst[881] = 8'b00010111;
inst[882] = 8'b00000110;
inst[883] = 8'b10010011;
inst[884] = 8'b11111100;
inst[885] = 8'b11010100;
inst[886] = 8'b00101110;
inst[887] = 8'b00100011;
inst[888] = 8'b00000000;
inst[889] = 8'b00100111;
inst[890] = 8'b00010111;
inst[891] = 8'b00010011;
inst[892] = 8'b11111010;
inst[893] = 8'b11000100;
inst[894] = 8'b00100110;
inst[895] = 8'b10000011;
inst[896] = 8'b00000000;
inst[897] = 8'b11100110;
inst[898] = 8'b10000111;
inst[899] = 8'b00110011;
inst[900] = 8'b11111011;
inst[901] = 8'b11000100;
inst[902] = 8'b00100110;
inst[903] = 8'b10000011;
inst[904] = 8'b00000000;
inst[905] = 8'b00100111;
inst[906] = 8'b10010111;
inst[907] = 8'b10010011;
inst[908] = 8'b00000000;
inst[909] = 8'b11110110;
inst[910] = 8'b10000111;
inst[911] = 8'b10110011;
inst[912] = 8'b00000000;
inst[913] = 8'b00000111;
inst[914] = 8'b10100111;
inst[915] = 8'b10000011;
inst[916] = 8'b00000000;
inst[917] = 8'b11110111;
inst[918] = 8'b00100000;
inst[919] = 8'b00100011;
inst[920] = 8'b11111101;
inst[921] = 8'b10000100;
inst[922] = 8'b00100111;
inst[923] = 8'b00000011;
inst[924] = 8'b11111100;
inst[925] = 8'b11000100;
inst[926] = 8'b00100111;
inst[927] = 8'b10000011;
inst[928] = 8'b11111100;
inst[929] = 8'b11110111;
inst[930] = 8'b01000000;
inst[931] = 8'b11100011;
inst[932] = 8'b00000000;
inst[933] = 8'b00000101;
inst[934] = 8'b10000001;
inst[935] = 8'b00010011;
inst[936] = 8'b00000000;
inst[937] = 8'b00000000;
inst[938] = 8'b00000000;
inst[939] = 8'b00010011;
inst[940] = 8'b11111010;
inst[941] = 8'b00000100;
inst[942] = 8'b00000001;
inst[943] = 8'b00010011;
inst[944] = 8'b00000101;
inst[945] = 8'b11000001;
inst[946] = 8'b00100100;
inst[947] = 8'b00000011;
inst[948] = 8'b00000101;
inst[949] = 8'b10000001;
inst[950] = 8'b00101001;
inst[951] = 8'b00000011;
inst[952] = 8'b00000101;
inst[953] = 8'b01000001;
inst[954] = 8'b00101001;
inst[955] = 8'b10000011;
inst[956] = 8'b00000101;
inst[957] = 8'b00000001;
inst[958] = 8'b00101010;
inst[959] = 8'b00000011;
inst[960] = 8'b00000100;
inst[961] = 8'b11000001;
inst[962] = 8'b00101010;
inst[963] = 8'b10000011;
inst[964] = 8'b00000100;
inst[965] = 8'b10000001;
inst[966] = 8'b00101011;
inst[967] = 8'b00000011;
inst[968] = 8'b00000100;
inst[969] = 8'b01000001;
inst[970] = 8'b00101011;
inst[971] = 8'b10000011;
inst[972] = 8'b00000110;
inst[973] = 8'b00000001;
inst[974] = 8'b00000001;
inst[975] = 8'b00010011;
inst[976] = 8'b00000000;
inst[977] = 8'b00000000;
inst[978] = 8'b10000000;
inst[979] = 8'b01100111;

inst[980] = 8'b11111101;
inst[981] = 8'b00000001;
inst[982] = 8'b00000001;
inst[983] = 8'b00010011;

inst[984] = 8'b00000010;
inst[985] = 8'b00010001;
inst[986] = 8'b00100110;
inst[987] = 8'b00100011;
inst[988] = 8'b00000010;
inst[989] = 8'b10000001;
inst[990] = 8'b00100100;
inst[991] = 8'b00100011;
inst[992] = 8'b00000011;
inst[993] = 8'b00000001;
inst[994] = 8'b00000100;
inst[995] = 8'b00010011;
inst[996] = 8'b11111100;
inst[997] = 8'b10100100;
inst[998] = 8'b00101110;
inst[999] = 8'b00100011;

inst[1000] = 8'b11111100;
inst[1001] = 8'b10110100;
inst[1002] = 8'b00101100;
inst[1003] = 8'b0_0100011;

inst[1004] = 8'b11111100;
inst[1005] = 8'b11000100;
inst[1006] = 8'b00101010;
inst[1007] = 8'b00100011;
inst[1008] = 8'b11111101;
inst[1009] = 8'b10000100;
inst[1010] = 8'b00100111;
inst[1011] = 8'b00000011;
inst[1012] = 8'b11111101;
inst[1013] = 8'b01000100;
inst[1014] = 8'b00100111;
inst[1015] = 8'b10000011;
// 0000011_01111_01110_101_10100_1100011
inst[1016] = 8'b0000011_0;
inst[1017] = 8'b1111_0111;
inst[1018] = 8'b0_100_1010;
inst[1019] = 8'b0_1100011;

inst[1020] = 8'b11111101;
inst[1021] = 8'b01000100;
inst[1022] = 8'b00100111;
inst[1023] = 8'b00000011;
inst[1024] = 8'b11111101;
inst[1025] = 8'b10000100;
inst[1026] = 8'b00100111;
inst[1027] = 8'b10000011;
//
inst[1028] = 8'b01000000;
inst[1029] = 8'b11110111;
inst[1030] = 8'b00110111;
inst[1031] = 8'b10110011;
inst[1032] = 8'b00000001;
inst[1033] = 8'b11110111;
inst[1034] = 8'b11010111;
inst[1035] = 8'b00010011;
inst[1036] = 8'b00000000;
inst[1037] = 8'b11110111;
inst[1038] = 8'b00000111;
inst[1039] = 8'b10110011;
//
inst[1040] = 8'b01000000;
inst[1041] = 8'b00010111;
inst[1042] = 8'b11000111;
inst[1043] = 8'b10010011;
inst[1044] = 8'b00000000;
inst[1045] = 8'b00000111;
inst[1046] = 8'b10000111;
inst[1047] = 8'b00010011;
inst[1048] = 8'b11111101;
inst[1049] = 8'b10000100;
inst[1050] = 8'b00100111;
inst[1051] = 8'b10000011;
inst[1052] = 8'b00000000;
inst[1053] = 8'b11100111;
inst[1054] = 8'b10000111;
inst[1055] = 8'b10110011;
inst[1056] = 8'b11111110;
inst[1057] = 8'b11110100;
inst[1058] = 8'b00100110;
inst[1059] = 8'b00100011;
inst[1060] = 8'b11111110;
inst[1061] = 8'b11000100;
inst[1062] = 8'b00100110;
inst[1063] = 8'b00000011;
inst[1064] = 8'b11111101;
inst[1065] = 8'b10000100;
inst[1066] = 8'b00100101;
inst[1067] = 8'b10000011;
inst[1068] = 8'b11111101;
inst[1069] = 8'b11000100;
inst[1070] = 8'b00100101;
inst[1071] = 8'b00000011;
inst[1072] = 8'b00000000;
inst[1073] = 8'b00000000;
inst[1074] = 8'b00000000;
inst[1075] = 8'b10010111;

inst[1076] = 8'b11111010;
inst[1077] = 8'b0100_0000;
inst[1078] = 8'b1_000_0000;
inst[1079] = 8'b1_1100111;

inst[1080] = 8'b11111110;
inst[1081] = 8'b11000100;
inst[1082] = 8'b00100111;
inst[1083] = 8'b10000011;
inst[1084] = 8'b00000000;
inst[1085] = 8'b00010111;
inst[1086] = 8'b10000111;
inst[1087] = 8'b10010011;
inst[1088] = 8'b11111101;
inst[1089] = 8'b01000100;
inst[1090] = 8'b00100110;
inst[1091] = 8'b00000011;
inst[1092] = 8'b00000000;
inst[1093] = 8'b00000111;
inst[1094] = 8'b10000101;
inst[1095] = 8'b10010011;
inst[1096] = 8'b11111101;
inst[1097] = 8'b11000100;
inst[1098] = 8'b00100101;
inst[1099] = 8'b00000011;
inst[1100] = 8'b00000000;
inst[1101] = 8'b00000000;
inst[1102] = 8'b00000000;
inst[1103] = 8'b10010111;

inst[1104] = 8'b11111000;
inst[1105] = 8'b1000_0000;
inst[1106] = 8'b1_000_0000;
inst[1107] = 8'b1_1100111;

inst[1108] = 8'b11111101;
inst[1109] = 8'b01000100;
inst[1110] = 8'b00100110;
inst[1111] = 8'b10000011;
inst[1112] = 8'b11111110;
inst[1113] = 8'b11000100;
inst[1114] = 8'b00100110;
inst[1115] = 8'b00000011;

inst[1116] = 8'b11111101;
inst[1117] = 8'b10000100;
inst[1118] = 8'b00100101;
inst[1119] = 8'b10000011;

inst[1120] = 8'b11111101;
inst[1121] = 8'b11000100;
inst[1122] = 8'b00100101;
inst[1123] = 8'b00000011;
inst[1124] = 8'b00000000;
inst[1125] = 8'b00000000;
inst[1126] = 8'b00000000;
inst[1127] = 8'b10010111;

inst[1128] = 8'b11000000;
inst[1129] = 8'b0100_0000;
inst[1130] = 8'b1_000_0000;
inst[1131] = 8'b1_1100111;

inst[1132] = 8'b00000000;
inst[1133] = 8'b00000000;
inst[1134] = 8'b00000000;
inst[1135] = 8'b00010011;
inst[1136] = 8'b00000010;
inst[1137] = 8'b11000001;
inst[1138] = 8'b00100000;
inst[1139] = 8'b10000011;
inst[1140] = 8'b00000010;
inst[1141] = 8'b10000001;
inst[1142] = 8'b00100100;
inst[1143] = 8'b00000011;
inst[1144] = 8'b00000011;
inst[1145] = 8'b00000001;
inst[1146] = 8'b00000001;
inst[1147] = 8'b00010011;



inst[1148] = 8'b00000000;
inst[1149] = 8'b00000000;
inst[1150] = 8'b10000000;
inst[1151] = 8'b01100111;

    end

        assign out_inst = (stall == 0) ? {inst[pc], inst[pc+1], inst[pc+2], inst[pc+3]} : 32'b0;     // Saída de instrução

endmodule
